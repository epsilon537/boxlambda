`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W6H08FuUtLHXyeAucIzI1L+gPAHwnrip7hASxzNigWkxfZQncSMesrxdaB80TYPhSCx0eI+WXFel
TnC/e6qXfoSiStzM8Gy+2eQxADDipEJa+SnIjUtjol9paVNi96VyPKgYNI1s0tVFmmWj5hslIHtQ
91MJSBrCAj36W5iwMgjUlBooPppdfd4RZiRYE+wd4iuxzj6KEpSziIky4b9b2L4SSq5WJOJ/8m6z
IRqoJs6EmpXIEdg6SQ+YH+cPn8hzjQZlcqpGHiT/tWylZkKGbEVWZatCx7Ql5criYPMiNaPLZBVp
yNQdPgBuvPNoldPNpYKnkoAMKfNJtHY0xlovAw==
`protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`protect key_block
NfROCirIvonjUtJ1t40P7suTZhmJtDmilKRn+YS3zVHzTo+dvf9Q10ChZAFtH7PF5VTrWX24SLkR
e113aS0TYkw07c2tFwheygy3HxPBw3NE17+EndrQ7RWbOREdS9B9+af7Z1dK2XVd9Rgw3W2St3qu
a6c9vBUUF7GjPWPFR269Na9tgc4aBem/qr+PPR2Hw9tiBg+JIZROJOP5cz2QRtOHIdO9ByBJNl/w
Ss2z6jhS1HxvgN/ynfNsF/BEUGMeUHu06s+qTRKxSCTuRkQK279M3pEbC/7RWR4FEZIelgtRf7jb
/AjCkeMOvxgtEnnWO7yRVY3eEs5zCFIxPsu0OQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Cb3/mlz4bynMtimgkD6Hh3lrCb00Wbs5Q8agiFkLpoRaDbMt8PkbC5/NloDIwUs5D40UqbcMDTGN
kMc9H1jQiQ==
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KOcvC3veuaVOntctiu8VVk4WNkasftk0Xx8k3gxQLpXZ0pgkGZiqHuPEy7BtXBdWLIE6RMd/yoHE
TK/J00lzlsIAPKp6FvAnF/UAaQsozTWG8fCEBQ/6qcU/X4n0QwQLPvSfUv5Yzl5GvU4rBwbusa5m
kdt1C/1JCGvcSX1vk3l7u+gh7sTXvL76Sgw6frbL0BlLsISoEXygQFAOLo+9WJWUXzpdl71xMmNk
HeX8UwHk74xijpUqpsDpFvxjb9tnmF1G+9xmSo6QKjqxP7EPKM0q5fD7W8yjKV60tOiwzIwFZJB9
APeb5jVs2E7Ha6hgsY2n9ZEUtsBN7H8fgJvUGA==
`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JTLBB5uJZDo5P5IaZjIFKoXHv9Dw9TWDvau8iucIZGHHE9VsnuZ8ccX+M+C+HDE8FXSpKap5ZMXm
dVHdluV+T8DPiXpQRxSkT2NeYWr/2Cr0ND8iuhoyninMdn6j2HhAq2nLVAWK1cfYwv2rJWGVxE//
8Km7yXCZeRIwtKsDhJH5LqH7BtUcLSK4DMcBWOonssKO2gv7XxqnBT1HZqqjq6a7pWDCDFa82ZLp
yK22+1iKCt71fuOx8wivtja3L8eTcvFXjgfaDK1PzIXjuYew51ePUTNFvO1boACB5797kZoHoF6W
cd2UGYEbeMto+0ofUStW8Y5kzoxEDv1MBQIQ5g==
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Xe9ujWvahFr6Su4L7FOehfmL8+qr88crtO3uC+oekJfb4Znwi2l0Z3UpQq/ATvySQnRWSdvEqhbx
S2YmU85Dsa+LoV1pG7xJMsvDgetPbnE1O7XvspqtDwfCYTbKxBGmH9YgyE0Ay7PY1u0c0gANDVCD
arGF/Oew465Qtb4mVFs=
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mzZqH4T64352/V1i+e35qTsnN0Pj3hG59HueGQ+HsD9jKMDXalCZjaPcLswYaeYnsdkydZbZz2G5
QCnE7Hk2qOK2ZdkkJOJOQxjIvlEAx4hhSYp7iKjVzEF0joI6GsTORMbnAZDcvcOGzjfUHtCHKNoU
tT8e41znIa4LJSTtkXz6wM+ZXC6gO3+IPwis0F+ZaqGVFISB58k2hR9Dp8PHDH2zP+XEtzCrGzlx
J3IXMNVRTiOX2JLPBWoCtDX7jP9OQ/BNpcxsrtNmV78XJMVvUF+ElTCeRDEjm4rEQT2xMFsA9EgE
SDy081GQX2PdeTu4PDG8AeudTQquzn1wnFhvqw==
`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BwRdOd8h4sw54DbfteCqdp7weg4tnvWKP1JcW+8HAZvVnr/GpOcZ7B48J+m7lc9SZZc6FgyalDZI
euKK4VdkYI82NN+nsJSE+pvJ3uZB1MVTKHFgFsJeNRijzmVY+AfF2Vx5XBOPBi+xNVpidva1u8Ef
8DhcHqoAbqU/G/Fqab8XYFcrA8CrXHMFebUgJPWoNGUjlqY6gRJs4aZgGdD2pRAw6dexa9tFd114
NB8uVG7emntmo8rdJD7VwAsXQ7VGHWMA+Ad7BDvn/uzd5qe4fHGYZ14r2CgOGl1oXDjXg9MmwdcR
EutrQTRUQL0f7cCqeGMEBNNWkTu1Z2sTLvde9g==
`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WJ0i+dcHLUwbjh/uig0T7InL4UIFP4K1ZVXCoG1SrAGEO3uFMyvx76ukHf2d4uKpmfq5BfchMYac
AuV4P4XGwHN4i1km170rVhqN1pSQlUEblgeev8ZCaIjf4toezAU3nar9qWM3cpb0G6uG09/MuPUX
vwiGmcTKGxpQqULKbs0=
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
US8vCyMOArwjJc9UtRkIy4tOfeLNVV2ldtEZCe/lgVmg90qQ8TuufT8FT6QkkDfdwZBdWOu4JeKy
+xI5E8skfyuseRcJ3TDSxOJmwCUxPz64UJej3YIPopRGCcD9Fi4DWmIogtiazET9qof5EuUFMnq/
Tbwv2QH+BK0JbsaN7ZEDBnliaoekkpurqOFjdn0I3EIT+exVNorzMkdBw50uE1skvUbHV45fBR4J
tWVWGwehPq/idT2SCUuq5dYV5E+yXDSFQMjsb2O+iNXRVuB67qPsGNcIXiXd6gZdFtRfjTbZ3MZ3
RsZTgOqUJBSn7wzkYcJ0MElzccVJA7kQlV+43g==
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 36624)
`protect data_block
2MEzrEtMczejxP4dVzxj+tI+2rbpiNPe4eGwFwrF7EwKL/FQDXf4w9iyE3PnBr4CtwXSeJ59jCrB
8BTHUeB69P/Z9IYGCl8IrLkp0xrUw8cSxE82c2o+FLxcw/iqbSNYKHMAWD8dTFBFh2M5N4Me5jQV
7Mnd94LMgS9cJZC6k/QxjYqP/rFWlme3d4b5+fLtp/kJlnJbhN5c3suLtpVUiqs+bfDteS6nGu70
mFMH6nzTo5qgwtm3/r4IaIpN6LYF16vBchTKKxmyiMvSfORbZInCZxNNnuQt4zR5ifItcrFrWo5R
EWfLJXiLxz1aJSB5K6zgjD9mWuGXePCRJFip9IAykIPf9WxRytECerFcGsVaf+uMPkQU/IwYzWf5
Pdxee8wBkMJEEO/o5LMaWokdaBAoiV6MkD6o3Mcmz2bbd/rwjrYE55pWneXFKik73UUAz5mKV9Nh
N84TK70nzfnsdN/XDaPyN1ruL5EoZVhMsjY5acTiVgZAgZeBRIkM2Z93Vz4DjmsM1tLVHHmD6yiD
4ZSeg9SDUwu0b9DJJZ+h01m3s9sxNKLRT8n0P2Zwz4dfWnEWSD3wY1WN12RkAmSp22uKfYT+vP6O
kL26JaTMarBAVHlIWzAb/gttCwAOycMdbJdUjlLysgkTkQZpNHi+idnl8SX7ofJ3h57Pi6e/o+Eg
MxaHBy0sdUHCfs+rd6eAtTC1cU5hR/gNtcoYaXSx4HXa0OkbLfOkZzfGSk6ue5dW9bZpZkjLVOJc
LOQgGnFPfFtyVCxvOGhk6kb3GobWqI1fM+D6jza06xFNNPtF9smI/uvPoukC9knctg/l9SiA89XU
BahVD2U9HykK3nBIDuYvz20J5iRCr8COd1bIuBiWo/FvYRWihM8wqE5vHifYYu9P3kjuRmO6/JsA
kdWbmQKCK0iJDcjNAl6qm5nz5ThDE5THGKe1n22pTn5IxfaU5FnKwVICQKl5tfXY2P3MNqcp72k4
f8VyU/5Yzw7jXyWpzvp6Y2CGNbLrGIgvmHDmatPAsCU6B9F2/T0vqT8M/e8C347w5lOj8bv0MSHP
ChtMY1XHLOg9y5ICuG2H7sL7lhWd9BeORtz6vpRnxviIhTQI1V6IVDnlo5GPmoSISp1cGcB5SceA
Os7OLODuBkkAwy/ianJvzN8XBZmZEW+MPMzHObXthLyG13m25gianGy7Wt8ZS8nvuxlhM/VQ5bRS
rcp99pBBFTUS77f4KZ4cWwcFNyBYXPPApLCfxmHR9BOkQ/LNN2GAO0WWg4t91sTlC9NdY24ueIsL
Wkt7Hs0bwCC0uwDBItFnhdQ2HEjgAZo5HZ12CvdZaFLZf2feuF5pfKcWduraBSXvqpGlyczHVMMt
wPBL99Wlj81cTrEXpj1Dn/Dm4UJ2+vnhfS5bPym3qdcBAo28/fjt2AeSCKzUh/kZjW6eU8YhzWKx
wTPDjMDHkvy1lv7mbzFxulVeGSTwDKO24wqslb13o92dpDmH6r7aGz03VfBEU7PM3OSFXPjnKb6A
QE1Vj+20sLL2LVpFiZcD0McsvYK34gD7hUT9wSfWTBS/sTQcLcMn5zgsNM3kGCOfVQMWOWg33Fi6
54UbymbZTVVwcTHqNLbF3T8zs9VvPgamI1gfQM7jUFD6x7CqBDkKl4GDpxclMpGXSm48+BAyY4dO
7G7Et+Cydxo/6hGiPbD3n03ootY47bGItkHNYPaZwXf4hpIA8xueFelfxeLEmtBhXpUlfbUichTi
k4pe33xfPxp1Yw1zSjUv475k5XIGKfWWQ7YdC02fL970moyTF+tMcmcDd1PJkPicnxUhx14k8SgJ
nZ3QRJ64im8Ci8wQS9KrevSD/fiSpL1nD5kheTLpXi8gFhX/UVQjxyaAvnSfUuoalw4OY4ZOzy+a
Qk9CTAeNeG28a8qAZ6zaeBbklUU25SlunWe56gSu8UTOaN8i1M6WI1AVjas+nxU8K3GqkfQxlXya
L9QKH68sJTBoJREiK3/IIOaz1a31mTu1zfQ1T5KySZuddURr4Tz53DDfxB2F4Rlp6c34l8uaK3Dq
k522Qm44+t26KeWVYlnfslObNcO6alg/FKTSUvOY6ayWsnhAyTsDb4eZ6g8Wxasr3q3TfcYX0arG
G3pJSBhYxW753qELykso4gTRTuaAFNy8mo1Q/8ZCreaeUgXCFd7NBkLYTKtcfP/157N9pnuqSarf
bQ2A/h3pnCpPTHnNrIrBE2SpYxEVo0TedbL1Nh6naN+GXr06Pp+QPYicyres9oHQwiD5Gl1YZhDE
mbC0d+N944q+3r1Bb7ix1W+r3gIkpe6G3ul8zJlSlbSepXiApJRdMrgJrnsK8NWekZsCvtMrTBV+
Yk8wQtXivd+NxASA9yoAZ/RY2LG7LAHEYUHaDe3v52eqPC1JMqMZzBb1NRLkA8/Gz0W4FWS9kGtQ
yPzy8NClOHClquAvDzOshHhCqWsKYOebIFZhzh84RoJGzKAFIdZjlBKRqsHr8n+UMAIooKIXEgHu
A/CczrdvTlGDL9OWneYRpczG76RrGDAyvkKDcmS6eDvmOmm7y4k8rouIbDqJMWB8RjqAiyjYxXpW
sRdD1DDXNar6p9qOPlWSkp+TIoiypjaEGMtutS9wMEfYivaMRla296oIZrzvImM4VAT+/WaZXpKr
x5y1kjI4EO25x9HmshYHjpCxVzhexrNbxumw3qQC+GLOtvCPRUcENjmqn7IJJbtT/d9+FmEcKe5j
Y2YSLW+rwdWTKAO+sulHc+0U67eCjJqGLBUoBbz+MPO8fIMobsuuT0o27MLBnvcG54FM7EpAIzow
AV7uTn3Av78630LAeXYXtyuyebxgF6wkrnpRqmjk1Sq+t7ukHrVKI+5OTfm7Anj7lgDI7Ooi0lGk
iL6nWeF4ZnVsbu/2nKckrULLfxqpOCTlUGRwIiqDRp8YJjF2LPfx26q88hczdOR6eY+Q5LsucAou
SHi1aLzLqe+8tijZMWLTKpOfehDJQU02cczzt7ug1UJvf9HhGYC57OTQj70+Uv1QkXRzMAoPGrL6
pOmtGVWRBFT4kzk4vtC9BJYCNMmWFwckrJLOP7R3Imv4t0Wk05z4zPdsLrLI3eqPqG546I76rYun
h2uCxQ1VEaCj9ygxmTxdudekLDOP1O/lhTIiF0qrWdTppf6XgWDZbt6YwQ6G/zMxTPIk+xgdzTEj
6rTSDkZrJgvzlUNrbMu/U1R4FI1BFUkG3MzVA/nJIWRIthC4MvIze1qcFhvh6apyVmGgcrzz7OF9
j7TkdS8Ml9a9zgqwl36KWMq9X2/DO8o1NBT6gc/gdUokVUMi7DB4bSWswUndFiCCjxM2qkaAkHmd
DuB7DhHLwu+j7H6j4pIP3l+QnnO8AgeWHUByt+xYhZg29MYXWpN5k8h6Fp/BuJBVSySViPfqvTo2
GE80vrIXjGtgC2qu+/6Qwyp74yKXhewc76a4eNFzw/S/0yi6lKnSBAAehtEtoYKxMU0012sGsdAI
TE6BghTudg22DpJKcNp426bbmZpUQ3wPosONA4wBeYwn3MLemvkKW5gjIVXsBVcXglFwXQewNHmx
6vYT4jeH4GZwpxzPPK0e7nw5+q2K46ePHZWViKkYlW1lMlGHxBa2KHO/+weIdlFFN5rU2ovfUz+K
unU6dKCzOQ+KEep/7QFNxGVPpHFpzrZt9mwQM8hN4e7kzi/UIrje+S1RMrzb7vyzkTfPzMcMWj55
9Gf3hsvU90LgUhMzWJOXxsRlFXSkrCUHb0lOAGB7q/6BFe6OyegDnfLtzh7/QkdSmS23HWt3k8De
QIKTnEPAlJYH+8yBuZ0ItXopyElB0hYBCYamoyYRbNDyJvKN9qrGYpc4smCh53uEq3kLFgdE1yER
RXmnVs9XUTTqCPc/+0+ZsGhmQ+9BjoZ2CgO1azCNWxfU3x9ovzzKt/Hybu4+eRda7jd5/Ra/Me/m
4tfrJ0xKhNw9rZWdWDZdiy3GtEm9bnk8g63zHVUD7xcgNY8VzT8QgTgnZaD3e4ZHZnZqSSNOT0gp
8SPGqqT95hIbmz3b++d3GNiroe7TfRZwFFXQE8L9ITHAb7dXZuBOyLQ78jbMwsCkuTwBHl6mHmna
JaGenoU7MVjg0iYBRMsQZi0Ept3iyRjzxUUnDJZVCEIqV5BHL/AYN/p6KU97mHKgVyytLTuk9bhf
8/eXvZtEiGjnZxeIaXFkZEe2Ml6WGG9HodFBkfsEpurkhGvgIJsEqOMsabCifP7/8kbr6FK344YQ
CMsZoukBq5gTCGB98Eu6LrGXOtwXyUuHSrAyseOFFYdqo0qa1UCuZ7ZJeJJKsdeMGlcE+ZTqAqEQ
5/jzV8hSBq61ElL4xRMWzQd3GT0P8oJ7ePzbKEDWAhvDOMEIaonU3uNq5UqkeKI3STal6eNhAVkq
o1Y6H/R6Jx8rTyqj7qVPNZMl3/zG0EcsiU7MsWTZjnogDMR/FOQPBFwLoW+xdPXkXzEfJpeGmCe9
e/Ma+LLQRPWgkdg041iOJ0pjMovlKjIh2EnzQ0muCHuPsKBJi7Hyr3k23mt+dlMl9/aWRYp2fuqe
D3NyBRmzgfW7crF+M5hfYL2eA3oNPfFRB1u2ZyiMIey8Kq9O5tkgOEkxTB0KmbUUtTgrL+Iyyjbp
M62xGOarnKjfqbFyICqhLkViQ5WgitkMp4ehtSnd53o3VEFPTDfa4VnRGkigAaiClvQoJe+OohfC
pGAfSJTZ/Q6ZVcdrPXDwzeEOu4ABKTUFRiDrGr2Dg2zGKhi+2rSBmV4QHK5sIa8nliFuAD0AD/dF
c5oMSal8OpZdrLY0oy5r498wsoZvMLgoKsF8KiDbeLOSAkFHCUfCViQiNyFQtm8v+p1TWEtIFhKx
lJQgeegBtvHH3zO9PAd0bDek/pEM0UL71XGdEDjKQm5JflxGrwKU8cLoMQsATeyUv+4xsaB2lIbL
xju0CCibDDjXanGCP6dBpP2gtCbVR936vav/mZkU1C/p2b2MrdCb0el4E24kdEWmX6kMsQY1+xHu
75uj8iiknLP4Ry/nhtHv0DCj12EhRTj8TR3LC2CEC70pvEfVKeaVlU3vWwXai56UEV1b0pycY6vt
dhT5CK+4p/0PhUAmO+HRwOGBl1AcPHXVJoZeQ4uMpt3oLfofMbdkRFzkY1/hEebjSwPHwGaNxxTO
Kv3Q0aLZOPQ07f+ov5JiS1XPTEkdODN1QRFfyxzbN2tPtd9kISlKkR77if5yTv56oSuesB5py4FV
Cwzzl0iuSu55YKbde60KQjXZQ06GAQlvsQGTV6u9jhaQi3vvEd7GkHbUQtgpReIL9ntY9ZcNKMCR
jCnhFTLHjMYiWFXZCVnYjSIbmwrwvMtQ3euCSWX0jgp9/ra01KNpsQyViprw4/ny8mEgGdBq1P6N
yOn3oN/TOzpw2gdvAdaskih9aZWcPQFT07+m8eSY32E8l5LrVn5wOyHZLZIvAlY02xG49mRKpK6u
hGmgGq00r0H8isygi7brl6xo8dOToHdmlm03ZwRfRuFZ6GgnmfG1P/CfwhzUQFlFnojKloJN/86f
DcKZhHZsOjstuCBki332yvPMs9yKhIiW8tzDedfmFctJxn2UEFE6M1qFu8HVzfSBjFHQAmMQ5Msh
frjFOipeWZr/P2WgLwXgrju82Ap3WujSJcefjVT2HD0wnFa+Zzb6H94Z0WjiUy54py6zUHvs6bIF
LbLwrs8Yx80cwaQXTMkgA4IbzoiLI/rB6ycbagf/tT85TZgJkNNVVCDzpm0q0NZkpmpD42nQWvTS
YMs3UxHz/YWrjlm54GpQ5BqIm8cMI1zJLwqZmxg951JU6ZSmI/xGonQCcxoUrKDk7CxDIvb2pwPr
0ToXzWEchkBaHda9t3oEUkHpk7UC7iti8B9LdHw5a8k/2wddX2SKz8D4IQYuHJTOwnUOcOoRyF9t
W1mrmoBDy10v8gcJYZ2hTbe2FknkJRCGkqIRYP8gqHQsa6/eU8ECniXwIunfRWSSXCv+hSsFW8ZN
9IgNONBkVxrxwgbQDWhFd6dQq8pGA3xT31jabJnrEa1fW/FEqvu4PfCD3ciG83X9Yb4D8N3P81CL
TKAt5qNwExSTgCC4y7rkrBd1b5zG/b+nhub+94uECxl8VkSdN3qwSU/OLRxwRG3ifDrNPgkSRy3C
Rw/dujDuwyeXH/Y3e7Ml/5aKdmkL4V+4tCZ43ew3WrdmLK+NVpr/3V2zTR4Pr+sT9V/iG5Je+IMi
WHB3bwJjBvQM58pG1kTuO93Rx6MccPxPKKcrOFQ5HP0s89HOIADHe3m6fCCx2E62o4UGIoS7hh4U
eh6ZbdFl914zE0EZXXY+gAc46r4ONDWHUCGczxVdkGwm1rJ1kTER9hEcFngnVssSdqjR7BW7XWSf
peNMCpFBjFV2T/GoPRlAuVFTDxUnMUCvrs/8z0bu5KJN8q+an7YBwZEyMf3IXSXwBIyslpc7yLhk
qI95lo9fUHuwljnRCABCLcZcy4ZAF8LC9goa5JZXeu2oMD4xERXGRi4CLsWb4yHHFZg3+xd2HobU
uPzN9IwfQfvLDVbqgoXSfgM7Ki6WX96P1uNctqKZBoH8x5isqZhVxa7YHkgQThZ0vOepG2g3XJ2r
qCKFks6+oDiffAKJmtjjn3kpCLdK139RbDHccNB57mebmslEI709vEZMMkokrAwY+rylbRlQZ/hb
qTRP/u/VxzgyskdRFvL4s3iBVsAfpvJ4lnHPpu1/nwF5Iuvs1HANoUlua6Sm8566w40NEKFqAa2d
6ZVgjhmJPhEO4s3/yfHZVygbmc6egLFBI967cn/4grqRnqw6UizDPOXfm2y6aduXnm+2B/37cXmj
O9pw//QXVkuKnQZVRSmF/H33JIuDOe225z//sKMELG7WvA1BShD5Z25Dh/vV40BKTSkuWkW6Cm/g
npavMXXDdkzJR0FxlQCbleZX2Lx21clvSq43W8jRHIPLEhgU/7PDiwMT0elRjLFGLiB/K3p3MAMb
u4t7x43mQ7NFiImedV8fpAX8REU7VFRP3IutLX+qCAxi0XzeulJdrQd7sMqGQh2q2l6kFEJhiLR8
ka8CMVfqoXK8tq+l0I/zts58b1ut9uwBuL4LK6Mog9FB12qWZTJ3Z3Vj6RUUeSSTaSy1kKH1uVoy
F9UYRfi9a5md2UyqyzFO1whRT4FdbuhicHPuGDrnjGMO2tDeu9E/EaDgMEYHRKuQLiiD2Nz1l1dh
PNWVJvkAgb1L3im+Oay8Lc6C0lZNHHk/XCDrxAMTJUSYOtqkUFou+Ba0D6IG6fGMx6QEh2L4GaDZ
39bJT8YyqDjWL9WMJ0/A+dT52GLtD17M4ayD3qm9M6Z3+eWZVhWxAuunZ7VVgJsjwJKo8SomrxR6
uT+f+YauqF6c9RXAFpdL/vGt1FBj9AK1F/dMuzf4ykXG3h+loWst3WwgDjiKjWG8HvjGvXAGfVSd
YbMhSZn1QgG5Xp5l8xrEirssj+X3EXWi9slM32753EQVOBV6iNX3sonI0Lp8pTmZC5IoXBDwKCtT
hw5BJSenC8Xp8qzULNDha10DEaE6BqjQFo/5ZLhjArTpPPbVJQA7nQdDbEFaqR8mtjt38kDtFgiy
7xVNtmRyzm/H/3IsHx/vi1wYj8ZhjoKKGCrHKXy+lyzWYhryxSKEAPtvyR0FgmPybVMOg0hxcJDc
al8LxiYU+wKY3acpPTQU8u6nghsv2xPM7cG6gBtMiUS++NwauDdJtuR71PmhzBNuDgkJSF9kFLNv
KStosCqEPgTr3Tv6K5EUbhwEeu7K2Si04C9ail/zjYezJ8AK70CzfwRT4XvAQba8VAd4icBzvEwY
6rq7Td/cEa7h1TE/ib4wpgUYTQS1lvmY/VVnwjXykqk6qHLdWhV1+fiEDjT8SpMwaSyuA2FGInLj
zkkY0oD/V947bnGQd4k61KzkZKAoNG+Nnre42yqKf0TlAgM9lw6kF+REy6kgyx9zFd+8HvRufPS3
jBIEzW7hJLM/Z5PYFS6AscxCRmLu7fRFlwU3/DCs/PYIBFpNSTchcZ3UIMDmT/88VudY+8hFW6lC
yl3n+PwA4lguJoYSowl8084xWBjcVW97xtLSAPgiDDvppPK20rw8j3STG0lmMzhAl35YDYnyrcoM
8Xd8xCtQh8RqJnsMnSVFO/iA4L2IXm1a1XMC9rDjD9vOZv6fXE0eYTQZDFbnTz4QaUQdGU8CFsT9
LgQW4TBCOuH0xZDNNoMCGUxUzOT+ix42xWtCmYtaAfxnYxUrMI1WpGNqMA2J1aaXks8WwdAbQlEd
Wi/Da9Cg4uNKhKBg5ki2mYD5ROLIKEL1aHV3U+ZOXY0ZsYOt4ds8wU4ZlZfjQ2cdCrTW5QHYxdYn
d2uzkOKgdgvnzsQCO5GKiSV5pUZnAG6NT8K/C+lDRK/EBETcTUfnBV6AvmldcruW0Sc7N6dsElcH
BHV96oKdwQjwy6PhVRKcjFdAm9wWJEGEp0uD0OlRdvMiulgODzoIgREpkQqiGymNOWHoFW5zit/y
djtpngyJLpaHea0yO8KMas1zQdAOBWPcXSL9Dr2a+8MirEWD6vhvD4Out6Uig0U3RJ+X/yJfnLqg
+LslUvkzNP62e8fDMg7w9P9EDrxN8SjvHF1JHqjOmCB2SGfD0kveJpem4uIyaLw1I30GwW53wtxO
k4QtghDIy12huojyy+LGDaZrWYUN6ZbBWZD4WFGN9eU2ugieLDpf/unT+5HdE7VqqbyRj+4Jyfkl
RKBYGbrkZhVrfxChRAG7rGmNNtKyNgfkixMLWOjX8dKsrgDuMXazukbopI7XStuxZcw1BqxOEkSr
l8VzR01w13/xOd5cbDwPkuDWo+lKQVvhNjChuu99vghq3jm+oFKIPvSEcN2rhQZ2pNm0cRHzFQnE
FHZlo6XJdq1+vZWjSu9xDu4jTEh/HJnE316mcs7ovXGVZRJwuCb7S33a4G9rDjt8JjiU+SsrW0ai
QUaBZL70Tz+T9G7OKctRI5dd7lWfQEY3s8hIWZwDugI6qO814x3GargdWg34dLJRNwQUuARDQbHl
BimBVnMkk3xXOcurNyxw8Hq18eICxwKd+brmD+V1xDrdWcIkz7JQ5K8GkvZOUZZUEzH4tJXEC30k
C32comVyAtqdupJILUeYEnma8tyRAedaYhAB875mg0cf5W7ozb1VrDvMvotATW99+IJZhDl2wk4u
kXPApM9SdI7sGBdRIJ0ID6VgREXYVXn9zH29OtjCjlhIcUJtc+FFLVEHS53Ry+LqP4B0UIW6prKF
0X8O8X9AlhTgWCKCxnLsLytQo91MgM7SUdj+bSPmeBd5y2XslVwjwpkKz1Ze9QKwaeWARaKx9edP
kVZVaAPEalmDYA6iT+25EWdcKNaH59leuVeM2NwIjJB+xqs/uPOMMxIzMOJs3nFhFz5wsU/G/jpX
l+i0yChzmcA4T04E0AlKF8Bt6WM9RgiiNNzJfesP2IyXcIgNr34DZ8Xu4FdggEtDbp0J3bu55VBw
CK6Rj2VSUlH66bJCGwWBqL5dHVqyaLw4vOIPPSCJh6Mla9KuuELT9D1Ju0JWtkCDQaM5DVyCIM6/
TuVxQ8ZtTEbG5kvjJ7lF+TmUSGDR0eZxcc4wZV/kuw/uz73/izD1Gh5/b3ABQdM1RncKghfZS3t5
irZIgFcOyes/uBq20gJ1Hk/hTKZMy2ZEB76c6xPBfjPV/pqXZBrjYFjAiDjoGOxQW8yl5Z5yUGFo
O1LlqXgbK1MVKOAcm81Li4CkhmeosZMH2dogR6LjdZV6VSPwm7NS1wsn92hbYPEVWZ8kKIoPrQIW
p00Vfk+AbUgoPuq1jZAwLxTsdYzu6j3tErqd2BGaBRQjN3wapkvgDfu4/YdXHWpz0a/mGSjmmXf0
7zPZ0nm+nNyT/BmH5xXORKgYgWXbhUNn8+gR1L86RnJ51RjAUUOCGvA0DtIOySlQY2nOUPrvZfcZ
ppQasCEKr7K9t9/xMVCryEiPhB/OckrqdcFUyLMiTTZrJ76OaKY31nAf+u/ljcFT9J8wNc9x6vOA
Gs+9zWDOe5PXvUKVE7bwm47qBBaxak2eLcWHlEHzSlpDEcuJLHhqx2ITYnst42+2jUWZq2wswGJb
Xqvk0x+WJwc/YKAHAGWgOGroC3XtYwPT9ikRpP8sYQ0f8cc3P+AwB8kn12B8kfQwxKsOdkeq26zm
Nj7imykp8reT0jqXoqLbNb+DklJiFfcrT9GcAoB6BA5i4YyBexLTGByu58iStHqfWt0D5tUwU6Zx
ixh8WQ2NMLqHYA0H/QiOwy81uwU2OVNsWLBeaQBGUtLFcNG1RfFB5TYp2w+medVtUeKTMaxNhXEu
16+zRsbaS9CwfiEMhlbPS4wg5zIaLRS3EySBRYe2agcgSDNSfGzMIZGl2g1cHc/X2EkuN55AQQ+i
40N9d1OJ9Vjor/K5mxahDLM+SgtupOJ+eeNN7v57yuREN6MQyb5Wl7vl6gnQYkYVVGzlwxmKODZ3
91Hy8e9kF9029CRuMPy3DXKnQipTSC5oD5Ryb+BMwKksCHCqrDkbe/5zgRiuNQVRQY1ReKoYE7Pt
U4mKcXZ45TJUNgp7X0mEi2vsgLH83eknqghx9bGMhB0CaMAd5vNwkXf/I/Q9QDLBMydxxn4OeLev
B50BsQUOyBK5WjuTXXRp/kk7m0lVLWoMiK6tjjnZn8mTtxbg514YfLb3o2oyuSaGW35WfvdZav/E
9hMzxdBgOPseB4LjIdrdQxdt4LIG4ruE9HQRx9TqN8kL9eqgksV65zPq5Wo8Oy+OmUhw6CgUazAM
9scYsABgISWi5F2nkvwASgX5Syqc2PNhmK5+agJES17o7ThLu6xo9z2G26X8TXfpAFUeKCbq05wi
x+N0Dle7ng2wlrZ+u2LnfexmJqmvfzhSljxAgQ12SNfQwK5Zr12bCUpRMIXKMCzlo2DkZCTmTcZK
bABdDBHxA5Lks5weWFAiiSmdx1DPqjsE6zSNgyI6u0n1m9EqwW/rgGZUjvJz30rSK5L+f3z3ISpk
6QJCOsAngzTscJbOTMOYOj+gO/PUCc6Dl10Xn+PFSflXqc6rCIiCku8kUGiD4aO3IS1hc1RbNMrM
8BKWKIY6ueTgpLNOtdlGLNkcn8vLFndsEX5B3lnLUYPLtNK3cHR89BdvWrC2DS7GbKi6WJ4TPga6
tJ9OUZ6UwL4D9OlCC0Nx6Du7973azXFSX6mG+B3RWEF+dAnomPCkHoZDAMCdQ0/xtUhYKVkDQxll
/CBC61/CA4VlVQ5F+xWPcn1bQI17zWK5nMty0MFNpA2WBtbeWGOx0RIaOu/nr4OGP1y+MUtHbSWH
kOb7DX0gCldQEExRSKgwZof2lkEUeC3P6PT2L/k9hD8YlBkMSJ7D8j1XpcvK3aRseYO+uo42U5LC
mXRSF//vhu0Y2H6gjnZSjhR90PFY52LIqRleA/FXFtuGZVWdlqZRX3255PoH0l0ZjKHHacLJ/lSa
B9EQespGScQoosQ9LufNZVRhwIyH2MlMvfkyoh7HPNzOvQDWWghcc3xV0d6s09eZc19B8D4ol8PR
+9DnzqHmirx+6VUfDzT3n/VVzbpY6CpjM7JG0K8fT1VZtnVrQ6jQUp0bEc1P0MmmikOTePH3+tLt
hBy+oF3puCipbYV7kgZTyRV1hZvjrr2lEcKhmfMnPCoIlZ7bLquXltNridcBVka+uyqpEJXxUlLv
Tmxnr77Oe0Iwkz6xt79bP9dtdKUTTn3+YyRvjjPg3hvJdwUPdjmwNRhWsJN9/eUi6Z89LvOSQqJR
hYJ6OunXjNpXJGwnzjyFpoL9eVQKzkkQBTBgKaDkUaRCi30MdmcKstrxwe1UZGSBOPec7aUQboP9
HuY/flhelE+CpcZfc4ciaMmQ9yGHReq4K+Da8u+SfPm9gW+KwmqIC2ITUneMOMntLl1j81Pp542c
7NSO6lEXOEhrBiaRFn1jk1UibeRHFprGBLI7SIuAzhijpRC9Ok7o1KmLQ8Sm2f8b/wRxy95BMu7h
mG4HA4JrSJkiUlK3PUO7fJqAKWluheK1W+psdpGxn9Zr1JtZs+T9GqvMbJ6uhbq6fQDzXNjrCubZ
MZ5KqUeFxmtHtnA2EIFa1iu2+nwDOWfVzUuuVD1+/loz7h/FtO/2/s16z2F6fNQQlwP7ll9Bv7Ww
Bkdk5xvrHqJuo+2F82DOyx8xZDVHBm0Bt2Xr1SyxSmyUAPc9VGDZrWV6t4HEbs5Ui4nb7E4o81cF
vuqgw5/rLNkBVkG1oP/+k/H7n+DpZR9vONkBNAd78DIuRJBS6McozzgbxgiNt8FYLJkMRKQHIeTS
/TQbiHLtDxZmtjbtLRxbVPVEFcOOJHKmMe5rW0mYplmbrywOFCCrRtIyAuEbZhVNEez3uKgjGQQp
ev2MSMSZKqSoBchgqEefZrVfKNxkW4q5ndQmk9F/w1WdNeCNiOUTF/CkmJbGpDK2HH/r+R53Ba3K
6ow3ywJvy3ELgUnWAYur/IzU2ZwBetv9Vsm6KCO+x9EHJN3LkBVTNMJi9uEwPtbXh9rT9HrZKVRz
SGfjohkWjoG44erNwZd4hlYjmJy4eIYrN4Qv9pDmNVHtlSi9zXlJ0XHjqTL+Acj9jm5NSjS3WjYD
rFVztrccfUk0wyTxsXFcMouoA0lS6RXJI7e6AsRP77PIupNGeC4Q4KU8doG0s3OH6E/zl2y1fp2q
nz7oWnYeREuuDqgLLhR/NhIPq9MGL//o1KpDMo8alB732xSl4aZ1+XjEtT38CcSQSXHlhBDKEUUf
BfYQ64CCfBhshO8wPwH3fxDLN51q5T2EJei9t4GPGQ3Kn1LJrMFRZ2A/zTnyEshn8ALZfPjgU90k
najG4Ble0oYyGKXAHtpN5sXYv5KP0/spt88dQS96bJhpzISqYa2ZI/ydpuRS11nr2n85KqEheBjl
Mh8QSRwcMW+VfAAzGyvcenyaZoX/11CF8aHetYywt4gQ1bOmE/QFBCyLRko8zLM3USasRsFoKWTi
Y+RVGgTTwzEP3Q95ufFSnjijzg3SjoUvOKMQxUzQMwvihSFYvZAIZmq1y5c5f5wskB9v5n4BD4jV
M1HxeBBrGRywH2p1maLC8SMW1WiIlMQ2AA0VED72nr5MAy7WqkkJGlpzIHEs8cmkSqJ/1T4wci0z
TcPXX6bJvb9pkvZe4v3EVwuxABy4W5wKR6tAXkZpqqxWZcb8JsCPGJ3ARK3yjR2hJUHEsOtpT6zA
cMRZMQ6NWxIdWCO4zNbNxhRLeZhnezQbbeAtAqD52ARt4WdnmX3icF/Rf1TcyfRkV24V6rSiKYgd
kQMyvJNsLgDiCmqGUJE1Y4Xlyz7NP5CWSVNI6GlqCr3lN0pQXYXubnix9qukD3t8v1+w7JpX+1UX
cNy4MD0zmFH9XiV3gxH4fp65zWt3NKLyd0Y62Wd+HS2VJt2nx+V2H/StT5FkY61q7C7bhVFpcHcW
2wbWrwnWpER46fdP0vxU3/77qfN7+uAdYnCeXyyiDZxkPsxHN++Wiwb/iD65RgK/rnCvR173z4qY
KBwZwJNzQ9QuksbJE3uw4xA37SHLogz0nYtyf/c5qq1CaSQ5qx+HTd3cylXkHIK4Gc8f67Fbyf2r
PyfcHSH9eB4vgXvf0isISsy718m8JQ3qJfQ1TnsT/TGt7l6GN5WP4cJRTVeRiLyXdmN6vk2d+ohL
1QUY51LVyTj6a8oWwmA/LBKB58IotHInKBCRRjzx1VWBPeIvzrUM/shR9/kpikV7V9+lHJtDsxod
/y8Q9UO6vnnXPebUI1+IecsWaxuA75sxh4Vp/kUonlvLD7I+LVlnj58eTD8AXShMze3Y3R2KbC/q
g6nmLesawYoJydR++5TDakV0vR+1GLe8RgmMaz9LbTEcIPHDipoBMt3lCFrjwBQNhhXpg+EGZoJi
8RMb/gPBexOiNzO54fPvNlhzklN4fsS/iI6a833dWnYqHMZoRSSDZJGBCKkFzl1fG70h8RJZyrY3
yXKKKRCvzIQqnWSLyIVO/+hvh2Jig19MlDUaxMnEY+X5cylIAiCQvDF9GYUTXpgeJXq+fgesnHVI
q0ZWEvSC216283AihzXNNjOWHN8Az9eQQ5tCl81Vdy7UyCn4xe7sgQXbmbINrvXHlRGQSJKACPvc
hf4NU/zSMrfK8QAUyBMCHZx2MblD6OUQ5R9KOoNJqIjcxrBL0yGyuIXzxiWrSzbfREPLzs3aAyeK
KGR9/vG0bVEqwyX9DYkWVNmYGxbU/vcv5X4UizJQThXwwbyO2k1Dhif7g3iUpTbqn8sSLgUVxBdF
qPuwbHPYipBx/LXfkvodO0cilojcOZIpV1nF67G5Qf9HQMykxJj8WC38sfB/KL7LJRvZUmmsvzW2
MOEYN5Fz0ULNcEDA1JkH+t18LEtHESyptKFKQ9/2z2nx7WsLic5FuOGhUUyFyftn1YKztvPlM/nG
+/ug+wNt1QKVdtXSK/84/uAG5FPlQ7t5RNqmnmzxDPnWJyOPiYzEA0cWd7mAm04j2VekBcjiJ4Te
B0+xqaxtoFkEusF84PwUyWlylI8jt7NfoWeKTvK4vJRNxQ5XCkV41e2IPcy5ePeWADLZqDTtiQlt
dFy3n6eADFbOU1bp7Z8VJ03Y7Jqx32u3Juw/iBOaVLA5WubDhYvGqkiRXIBdXzc+K4dEzgQMw8U1
vDww0SvlNBCwO8n+7uTEqgk/ehC41x71qj3Jwd8RidlLAisNi1aQhzznK6eo1DCXikL47u5WkTuk
3oxrHvfoDkDo2EqUbBBzXaDcUfWrKC9NJ3yrAk50MNOZwgl1W/yr+yFETqpbzuWTZOVHiicNqVnb
uBrCYYZ+TZupdfrbrOT3zhsi/feNr3mTfFsbBTSenoNyYlpc1cPBuQ1D7bu1OJqYXCrmdbLn37E6
9ctmZe0xxXryCqE4sFJtLii1pqccRui3Z2R63pXSoqtUnJTGY3tyVWRUcYBidNryYEwbKIkpD+c0
zZojBVS1EfjrcmYFo8t+y7HHSpHlCsLoBxm6zm2/t8y2Fd0sWRBcnPi7tAh6lQSDasZ9yaimKJcg
6yScn6kn4pP/3+dxJbOTd/Yb1GW3FLMlPDnLWAQs2ktPNLi/dTrrOPpC2mDrGYnijXEfhimBRToM
qrRMr3Qsf6dMwU/SYBJP0zYkbMr96Fsq5aXgq5+yz78jamhjgf4SlWEn3t+sadfsXen0qaQE3/mL
f7z01Jgcyh/QVxq1vQd14vMDdW6z5JroIM2Hm0yfgygQWBJnc8IKkvmejOiY7fx/qtGALR1jzokO
+zF9PvXjZVBGhUKlwxX4Jn3Pr26Nk9mNPkjn7ztrh+V811xLAlOgVp1azerHzMO1fBGbu7snwRNP
XymMvB2KWLuKJI8Xr4Ohra9TDQx8z1y8/MpEOEwBSM9YqIfwJhf83anNKjxnxXyWWhY1XnGfgxYv
QwBq6lpVkQJpXBCaeYP98pXvv0hNy+HtuAodYjKM0EFWQ/iOQ4jPd2JWmtGnKS+FnZpRkTU8n7l9
kGlA6KzSWDXqphyw5SNLXOkrVzDRCdLmsLk1gkFwM8Dg0jjWzgo+9i4t1fOJFfYgzaMFq7xpKSkI
CLMRoQlpZp9FinY78lEfL8s7q0cqMtImdgAQ8tEfHLnb0aJrA9b5KCoXIcOlVQPwprtANqSfnfbP
6udk59VjOEz7t7r0BHjKnpXWBRE35CscDCmG2WR2AeZpmOW3UOcnJ3b0Py+1N4DWrIirIIAOrBZN
aFCsyqiee5fToDuhyH6sEZ77Gk4A0d6k++Gsm/+JuKnWEJ9BQfcfZ3ICmSWSo+3B3rCijPb5ossR
NMWXpW7zT+A0/9xjg/uzunx8SeSxY0Vy/RQD28isEfnZVOg8k063R8NcoTSKXC8wxpq03nyWxQlD
ut2MyYQ4nvHUgH8VjZNtjWt2cLJgziWnggNIAoSFU7rKrfBQlz6cb1x73liSeAKe29pniG/Tzgh1
/rVLR8KmVVhj37y6s7QIYYW1yRpd4prm8gtzLAfzg1sRwPlWAVXbZSBwHyxdS5S1Guempt3q198o
1nH6x86crXrsyFZ2/zWiybrYc4i45f9EQOtAatIGeSBkTc3qh9MP1+kq08t21O55z33HQnNJ8Osz
EX0mSjd8tbl0zCkzZZrjTfhwftPE1f8Tpb84jyLa0rhGpU95Zlp2Cx1YJn/aBrG7vHcX8TIP5cx7
KwV/N55GZ1ASDhk+SI1tZ8/iZ64jidzJ1ePA1RZESEWbEov3LZa0kt9k7mMCmsRYu+pcjFJT6ouQ
lam5vaKHpgGdWYj6oxR7StklvrC4j4b4/d+OsiTadsSDwl8crNQmTav6JBsPMEspqBmp70MHrhq2
HbZHqr9PN8Mej96XCTVSzlVCA737de7x0gaf+k2a1s3h/QIkz7wpX9LRTy43YG/0NoHsUIHwNHVK
StQDIHC2XJAidu1GFH4ycqQoRCYOo5JC6EJiTSahI3wMRdBJ1VcpqtLpXjZ6DJnOI0QiVqcfhcJr
zX/BZdaCd18AnXYulIFdxgHSbfYdTtEX22y1xm3ZUEzPo2kDKYBRsuILj/R+fRkGpgSLJWsR5wAQ
9pvZxPj63sNAP5piaq+djeAry6qchep3c+tJTxWHvslpadWEAcyUNzHQy4wiyQFgmI2g9rGZKoKH
W8BywjzqZHTe/qQV9tKFUgDNZckzyDyzsOmz6KCzyUHtrLdLEHumSsco+7uEmyFAIGe/cYof8rje
siaqFIQ2yR24ivLsrbF3goGAPQhFRZHS8CrOY6W0z1MJPAc6zTK5TKarsSL8Fek1Tgx0WLqrwAvo
xsapzETVpJqGPMVtvX7teoxTU/RSRCdeIhn8OIuhlrJrDeL5/9dGFd6pE258N8Zg/kWFE4OWaGGp
LpGq18iDhVEfHBn/eFQly6XMEIwuW1UuQbL9vYKERprd87TmcyD8MTROpcaslL/cxMl8y6C48ZtK
AgZ0/XOe+O9GoKLK0Ro23RjoTXmz6ADGMhNIv426dnCCpWICZjCW/S5+rPw4V0ZBqbyQKSYCAk8C
7C3oUy4Rer/y54lQjWyOJdCPSvP2eupkSf9nXM9tSLdRwLbDMxaGSaH2ri0W6Bop0Nz6pkQNQq3R
97nmSt/WsD75ARREQEqndwd8QiXo/zuX/6vPTjWRWbCyF6gPu4ZfTjf88oSvNLRO3QLti9V5M1hz
Vn4Vh+YghCOfu6Px3h9NuQlf0w3mnFlUVH/Nxuk1S+UzT1esdaXP89g2AzLcJOJjAizzlI6CMMBo
WcK92XVn/LqDhWKTbZdpjZX0LipZr93UyhUujYFLyZEeIHZZT/jHZJkV3+ARPflPkjIXDtifsP7w
YwnM7hrW0lGvVPx688VHCb1YwAB51OL8sL7EHKtFFf8OiRNxuM3CLkJO2J5OyaYI0s01KKPTntMT
VPTJLvyrekay0LIAB5Ri16h9N2Jx7LcJ0vKQbFPunxQwPy5zDP2AVP4HhGWp9DA6kRpXs0n3A+F4
WlzVo1IOGVoZ5Kdg5T1QQSPI85H/buiBk/ukJkfep4P9nofX5V6CR/yhTT6HdmIoGRVQjL4Zl9r5
vK/VK1berWQSf5/UZvkBwzvbSFQq3AIdCIoQbtPBy5vlvu9J2DmJ+5mZdjO5ddfN0gQngpEJzvSz
xCojPOKbThOvqC6wjf7iorq/70tyG0hjj/jn5dvRagaA6/smEuA2R2tHXrS56TjsZ9nscX/CJd0d
9ynAgS3O7WDRIouUsqxRPQvY+4JFEg9K0tBADuslUP5aHESa/uh1ZcJHRzvOGeV8NIOfB3jaQICm
p3rpjfnZ56ivXI+Ivg/ZEU24WW4gHgFXfoF4Zes7SvpthP9KZ9xxzPdHrR1d/82Vu4CsJznXE9gQ
D1lR5nHdEtE2FO2sUHlXsLsc8+2tSPtyppnj/slLqsE4Inoy7gzVgGNfhMFoeAe/SXTvuzK/p1su
3Mt0v1p3z664qhbABtwTnzh/Bg2caSdUZ+PLnesuVA01GwuD1FYkHRePCde/HmIVZy+didh9nXx6
HuenSyFebBMkqGGwydLaUJJB2lxVlu6Vcn6qrW1VI0nojurb1suoHbYO+qf1pUsyjKULIT3QtBk3
ge8siHL5tiMqLVY4aQcuFqt1uW8Y+ZLSj9PqQUFpYCHIk6bLcWXV09pnnyeY59vFWwoSlDuBlWhm
zUSvff2W4me+2RbJpB6/u6B4IIPhOuJybphAZUZ8r6ciMUAEjCxuUYH9P2zWdVh3jIARwp80a/VH
sQxkZchnODWqMFB+q3XlYFIi3Sf4kLISRhWBTn2CPG+kZxU8Lu6A4idPJ8HzUf27yWJCEFeceCRc
1STg0w5ZIjyocR72W0GAX5XLik6tEkjURyndDD5ffsCrjVieHkTp5e0WhZRiqRVGyvAq9XC38RP3
M8VToGQ7M3rASTzCwVkqd/AyhoToHWm83YqrtiCyRNaEK3E/OVJYOsb3GEZi0GiQqV3LXD9/GeIK
f6ei49lQhUeSngIMqebCxEYBKfFfG7gaSJHhtrVdNGVo7oxuJJOtq3cIWRrQkhUQO4TUrNEd9M6w
6pcsCOqn1qCoE+3A04MydW6OFud2UdoUT0MMHdSd1iWs4VE9HldLZfXxGsWU+a5tyhDUzCUy5Rtp
RUswe9FwMqi888oquU3TYW+zcyO4SpiMAm+C1bzRC3ti7gdZnH/R9dFi+QdCZVNrvTbGavO8WeSy
Yi24ZuG8CS2YAPyPCgt3klOfjx1CAm0MpaWf/FxOQwDxLZTiexgQRGnuJl/UKNZ5KpGVv8vneTJq
YNdINi0d24pPMJJp9h1XOm2lugq4j6BO9uK2giQjEh78GRYSKePBS4lWfaCBhUxt2ztbfvJkKCaM
ysxcZc1GHOfm5fvhLQLr3dNCMf4a7JXzNC7wfp/GkZIzqZzn+CInkgEHVhcMB6ijDShGm+TR3X9d
Qj5KaxlDgvm9GReTkPUOK0nXlsigM453ELylnWrsFTOjBD6Nj5wsRF3HZxADn+5+NV0kip3RlYJS
0xwP0KhO3qvNkJU1hycNz8OCpRa7X3COLj73ZimfEVXRC7NFsMOxP8u4Tt/yLILVzxtHpqPdMzFm
OGVuBoNhuan5iFmhgqcdQ6jxtucA/ExVZYBdtbMaUw+23023QdLjER2G/rBpQILuOwm7bTg4lAe1
qOYYUx2wkgLcAzZF0+3ftLI7lsZ3lEmcLoa6Sdn4Nw92WlrBK9LgQ+6Zh0n1i2HbTtnC3tiMbDuI
mFx4uIYaqculLDtsauJ7k/7xIKHe9Fleky7FGXa9hwyTRQTo+JI+QJj46LmokBOnad9FWnM+gjP5
65HIIwFTz3zt6vqsV0E48QZn1YAmakuDOXTUy5xFQ5UkITD5ox8iYWfWZCiyoUtj20YgbLYj2eaS
QtZZ815Rv6BamuzCQcnuaynYG1JbzM560s7V2jXYlXme2407Xsi39reiX2hj5IeoajH2YSL7Rpfk
VC4V9asMopZLRXn474YiRcTtXDcjBvd1StiVTrMx+C/U6SEzS6K6liwiMNTwI+9KcldU+c3fsSrB
lfeQL+E4grwbSu9lDs6oTLAK7x3JPvNI8FQFE1VUOY72axULFQiStsHRhQrt6PWGCzBHvaStOuIE
5c3oZEqFNpGAcyQCYZrUi4rhB9ZtsDOwReUujW6hGMZiHZ72edyPcxvmfXz0LsFvtL/J31HVHKdP
GRJT2mcPv6xFcpbl9Mbdp3Xlynh8dsf4OMPWyzhmKyirF9hbvvHvMchT9ubPctWfaXrRA8nHAVD3
ia7bmFWz3/lYz6pLkGThEn0kEKQsfKNdBLVOWV4aqctTu7rIlK5EEN2a6ypJ6lwsaoWTLRs5V7z7
xD9CLrgeqL0jk3e3NKg0IU+n3BeVLjlwOFGWdlxL3Hpg2qQ/O1jdzC9ZcEc/CZqkSHjXEPZuBPnz
pROP1DJ3jGs/hJWUfnI17D4mkmP7nYKc3t39XINVErQmCvmCmxl96H1rA4XpRfLbHctW0D5D4eJI
deStY7LKFbhYLDNTHKAoU1uKrluBe0w1EUq7hBInheFOkr45MVQYgqJtOfSaRTkPkcb7IrL3+mAp
4IRMlJzokqKv2/hhGzYxpjBMjSdq6acRsbKnMTPp+5PcC9o1gqYGzoGZ2n3mHTo9i1o/+tM15DHM
Gqv2V1c3ytv/qToz13ptyWSm5oePzGlNH9M3YaFPx9/awiIhhDn8KGj4wfo9KJIOqgXI/cZrznma
dWw8Lc11stxn4TTfOoAzALuqi1AJ1mKF7fvvSi/xVvfxEXREuyS/zXDng8YFbn1dGcozYYlzLuDe
zsFcQ6JiefhUoHTAOgOp+GeedsYbs7/94SPp5+LD6vYoUfDtVyq93RXUjhxESu1hKFxWAbFQgQcC
EYk6N4IwiO0abuPkBnPkdb174MhbpsgJfzpvRQSTowYKvJA6IlBeEBRJycDrULaRtFxFuWssdofr
qcAM/dBU2yfRDF0nauaqaFQJ/ZIBMfNiMYbx5hokFiXcpF4OB9pnQT2RFc9G2ka4NZwh0ihxMesJ
vNdEzdH1FujG6tS02+WuyYh20LV3aiUMa2sVGaE8e2hyuo+oj3SguUENHNrQErX7RO072XiTSOr4
/7ZsUJD8afegdS0ZBLWmlKFYE5FWDsex4SXRNp3j1Z45ASsL9oQhL+APTvg1oH+4LJDR5VVavbHR
UOm5yI/iRxo2UsAGmiVBeGviG/HXecueTc4z1O3XLMaAJX4TqVWVQXAfzyQqjIqcSKVsFz7VWNMI
0pS3PBkhnCCNW1dBTyr6nayqPEnan5O1GQgAGFRIafpBwQabBjXepnbJVEaDsOJymz3uej4X9BDU
r3xFijJ9npEAkCkRmHexGXQhOljSCDOUK93dJire7S9fmNgQubphce1c6S26mdr6xz64VVxCIZCh
WBmPSehOnXK1LXhkz98GEilWcfHwY2N+e720Vlhm5rkhmXNlcYIix5AbtSK15Y9Gggo7FGSvt114
nzX4vNKdlWhHVrCfUohVeoeL6bIlxYPBPh4pWcMdvTt0Uhyv0NsFOeJrL3vtolzB4PKb1dPW4C1W
RBvtJPOvrAH0LJ5YW9J3HmkJzkOnYsxXTwmBbPXoqOB4SC+44tyQI3e86+VThFXCpMD6E1/t6GQT
b+zj7z4KEIeDMZoZcakQuJxOPG6dfj5mwXApv0M9rYRFURPKoHuLIBoGDvrK3vQxnfkPeBuxNlL2
bOcAw2NR/lub2kRS9I6Wx9f7XKiiNEnUanyML9m7fJqmzLiZG8Iqt20C0l+xnaHPF/GFMc/VpVwA
p9iCmSK+TGhZdsgiblDs0f93dvycHtlQ5ndb07f++eJRKNu9bbUJqU8qTpOPUZiGx0MennPosVKl
Gnh3SQ31jRH9YlssdRLnvwvZIMKtVyM9hsZpugS6f+Pzb2ceOfbev4MeHIEgPxTvxCBhIgTTxBIy
4aNSb7piUVfroIgt9nDO7mty8VSLQzGiE7uQZADbf0mECzhA4/EaB6TBy9M0OQkM1eXDbD4wyDUS
SEoILJ64Za4euy/43S8toPz8BG04HZeL9eCh2SxlJJ0tWORNvbM/FWO1FihZy+b5deE9gNEA/yGv
JuuU8sq4GRjxhOd8eC6r+ZD9jhOaUnOlzO182/f/gAIweeHqeb4Hl605fHPMxhtNBXYWikv1LjLF
jec3tnEM3nAx1Drc3awo6q7vsM3MOxbji/cPKGFE9h7iXYcOx1XrlAQrshd9Q26r7ha7Wlt6eU6n
uVo2ARfgiTKWfadcgncGoxQzrykOcJLQOKzF8hod8B3+BIGUvfu1JjzeRLRziCI2IWV6aEuRTj19
eziSHTvCYbdP3RUKm9hxZj5IlGc+gOsxHC12CNHKV/t/eoZPOLftgYYbsz1rxxaWo6L91uGJlV3b
CLRsMZ5965IM3cQ3aUUFCBEUT95G1yvMsQQ4AIJZh9uK1EqMfqwcBQMKHJ7czoJaY2pNCd3FKngu
xApoMPTOBAimr2DsniG+XW2bIYtdNtZerFH7ZCQ/J5qtpk+ftCTLJ5IbWuD1q3fwmG+MFbggQTAh
ElKzt4BvTWmVjFUCSvubuQoNYwxDvtUfBFWOROlGlffb2w55zPv/5XhrGUnPB6GjX7RbhnRtr8Jj
ZhJrHM1i+kjPzlCeepB9JQ/UnAuqv8y9rKogXHaUEKnqW+Lm/NM8cpOhfoX9cEYb3t17cvYqM0PO
7BQfXraGE2QMTgOvbSVKNVePvCVjkRgTi+ZTz8B+9jR06gjWEFD9rcDf+r93kHo51aAA4B7f16+u
S4ZAvEljitcfTuVuidaCzo2ZWw+cp3f6O8OIF+OEC7qUah7VfaXGFyhY7qXiXd2/vicTJU4Cn0n3
2exxCts5gwf+WTT8zpPEqdkC8QJRqLA5hzPq3v9wS+75Ktyi9WTHh0LQkk4fySUBFG32H1rXiRde
3lL4Onm0q5XULPow0WFmq7jcoghSXcjoz1H6Dlzb4+SWCK/lG/YEYjRxxHtOdu+MyjSohhTBWuNX
hlgzKMaJNeHh2xvC9pyB17qh4g4N4IuesFKxK6ryc5/07xGGpMEhC+d4T+n7Pgt1d2M1xS3ihyyK
ZDHKOStln4zKQGAAOlGxzY9aRlZKzYYaYHSX3ZmQ7wuYejwLwpiU9uzvqMD7q3A00VoMUQvtbwzw
W7u6ZvzWFjLTGlUo/+Nk31xUWWuYWasgi5DLPLXlyPPS3+i+Zi0FsC4vRkE7MtKniMQl8Nl73gBs
E7LpugsvJBd9lbfKj8aawKc4fbDeWhOPyr94X9rrrv4o75wwc5FyB+2wmtDW/pd/WnogePgRFTfO
IlK5QV73p6+X3KKkVFu5EgDFJ4O/aeieLqfNVkAQGQAdzkN1BVoyxBVMnw3RppnYS2JshYB+5d3h
1LH1Iz3iDFbzUxfvrUCR5CNpaoFYQWlRWtrPFk7uvgbscZYQKIt4HbQj/T02TLALqpsKJFsIj0Mx
7btzoghkygfTHuegV9zywePHhtAgmpa2JE5ewYYAejt6J/TiM1safBt8CtMpdU7FMPiW9Tt+8wbR
DP4a7TU6udxbqOIvztoR0sTRa/adoEt2WlBXiSRRoWNYCocQQiLTxpJteoWuk0zilHMAYg6YW8Kq
BenOdW4jCwzOpzMfolFFbTAtX+zvfR1Wkv8iBsQHdYC+3rRto3DBVugDvAvxqdFFuiZwKCQfz5ow
twcAQswrwpVmXIQoW5AjqFet1UHB2YX+2xhlkznRE61uIWp31KdnrZ8Ulz5zbeJpP+mivtO+qyEp
LkUPgdrIakW88UX8P98S2FFhpcH66hAywmiOqLmMvPRNxL9grJ9TBrfrOfnEQkPYzcOXiUTEb8QU
w5zMrbpCZKg0BQlx3N/OzjtQ0IwEHNZcpwPROwjbzQGaPjeZMwKJk4VUjwQGDLJYfygUPiJxWOJu
zqPiM8VygiUP26vVUMI3AZH06Uj4FL1UP/sTUQdR57fYTYCt6SwRuWgmOyHOUB4X+wjjuRCWnk8B
hjCiwcKmqjHwBT/k8tBMm9dIVRvmw4cD5PgpCyc90sIckaA4bATtgeXR8UoQCJj7CoY2h3lyRpIo
SGX28B+CPMtal0A9Teq1gMntkYbxe3sPQ5FR/8mie3uXJj423f+d/r5JMcEWxOHYF6w3ng5olYPh
S7GUQghWCxWOvAjrIn+hRpIty0Aavookm/DWXdT9njY1+g9vEw5q4lWeix6DnCBukg+bMPynjnKs
tbeA3tVHX0cHyk7i7vg8/pBs2k5D14DymvoWKXwGynYAxwNiZG2A59ZyuIzfqDPFt6819LoogI6a
ruiZVKBQjotZX2nkHPs1Wwt/6+QL3bqptTtPE9O2hz+PKjMBc+6oBPNQvgrxECjgk8P7W9F6kZNK
HhrRTfwdfVzSMAQswnK6bV79+1eVRIxivhnacQZxVLvslXjLwIZjzOdFzgdtLoAkqzWDurrVHwgr
aE7Dt5rEIVLG9Lp9aqEZmKlrR57c4lNuU83LY1zzz6//cO6rnIWIo/hXteCufw43zFJgYTl0/Ym2
+X03wpQlVPdLyEzSeFaJ5hIUaS7oTJvnqw965uW2XWjbA6p/zgR4ng1zwcU8jHHemH/8RRc3dAZL
zRiMEc7hZMmg8+maEF9CUD87Ds14HLPpcxMa913pgC1pTv3d5blK4X/kfp/PQ/TPYrxuKEmOBBND
lD1++2NcnZ3H9KecDT1oqOxqScqD58oI4QEM415Qi3SqqbtTwVqmD9dmxLvI6SWo3DQVJL7lQg6G
YrGD4hWowSaxEAFY8LUVgFik5sFgEYzBIFprhRrEyULkjP8Gnq7NO02vCXY2aNT9Z/BdXCV54vYJ
esr3uff+lL6mrDt7wSZEEqXvc/93xDba4Z73G/3/nBfGaFFT7G6oNQLkTHCC1z6vlrwJi4lDVdrO
JYpgpgqa9GFD5XLEJ9+X+GxsmjXP+qnGddwzX/wWMln3tvhirnpBvJRYs6BVHzRdperxMQjfMVGB
9in0o1HHDu+vXMBkgWNOoIX/QlxVeuEsCMlibrZ8dTLskFm/z9qqm9Y9x/dMcT5tfwRsO5U1wvA1
SaakOkYEss48vtJDFyAzSe8jjVfXwdxqn6h2zh9X2iatU7AqkTt1T3pcvcS6/ekGpG68YWYVT26l
QZlUNUC7oYcxB6gcghEU+0qzC6uplWKzruBRVTSOhbOdTor8qUDR2Ol04Wxas1BOayVoaX+Z54IF
bqz3uVsO+oLElu0DSFMLGSbbjzfvM7pLdBop8IZBwZ0KaMie8XeyT/ixUB6V6GEf4rA3jY8v4Zu0
dBbBGr30ZjpJpPZu3ERjfSBeWbUAVRSAW3YS4zqdEHvdcqfuyXg1PE0jzOQZO/NcCOyrWqgQWV3Z
2SXQdNeyLVdvNWNqmnXW6mRcq5WO3Uk41Zhvy5iQrFtJw2qb1oe7geR8qOEZKrnb7wLZha8rzhri
3L4aDIEG5budrMfSXXINpoeCXJmxRanFpPxzzxKs1qZoIAQbd2LjvvhfCYLID5TC780ciRf8Gydx
y8oOAlNusdl9PyC7R2j208iRiHEEYJe3TcQ4CQH+fznLEFrXdXDk8Zzq0vHWxwroo5UQevYMATtT
yUU15iiiBwJQoIDVzJF4g+8JNIVNjkEMJEd7ZZLKRhpIiVP1xmwlc/CZNHhA0BWRr68h76jslHvP
xCsktnJOgdNWNH2moxoEkTCAUmaBlKP06GSQ0gVS0Mk37ZHcTpHN1n+R8RaNx83C4wMHCyPiMoYV
BNmI8x9RrqaN88TiZwROsZ8Egi8AsGuBPxbkW3f2KVhSGGsrBPUbNqbwWHzdOTQynl75NMuHsi53
w7+TFVRmjZViwSolkcqg7i2Q6aaAFzBzuaLIMhcrQwBid74Z8Qub6KcjIDOPbIR8V4isiTxA2P0E
ZvTJSBSTzH6Mje2Fb4PQGC37sqVb9M8qQgY+e1T0VvnWWBk54mKNlmvCRRC0zmAJxgS53/64gNRm
gzhB9cd1XnWtq7CXfROnnimcdkisz7a4JA0aWbM6tO6Chqd2UupvNEufNoQsP1q3Muc38C176D6/
aDxiBfWaUjFQ9rarm3Mc/UkRNRqLY4vZ74aiyYZ4rJw+bV4r6u0AMD3GlREG/c53deBen0o3XY9Y
1hW2j4H5A/I8lpCkEDdqUiQXzVCq1Sx+pzz6WAgywNjjLLIsGn47fiAYdBHMF+jiLqQel+bx1yNo
XarzaSqCrQxGwh+lfzg99QVhWp1jcd0kC+BDthuyc9mQ0rvCWMpttU0wzbas9CzknJ7OHe6TnXn0
63iA4RARVuVq7dTYvjghxmKIZA21GEsVCJO+vijj41/54hPAcl3xFCO7oVci6yVXwlFmnAVzZ+Yw
JAUe4136NvRMN+nqG4E9WjThqMZPvL4HbjD/hx2wn1yTHRt1+RlGATfxulyYxKn+fZhW7MlU11PX
7pIqUAhMeCHQpCQSyJHmWYvMrAgc75glBLd5DimO7Q4fNaB1i5St8wJ6Xw6JCH/YbR/ghU6JuFUk
3rW7hx5QdDd1BYohM9kErENKKwDj4abgns8QdXPUR/BrT9ZVLtsnprwHIYRg1+K0pnwkMyHBlM28
HAzSdM7jTucGUdurhETsvBq5FfNVSf1MsHkaC+LSOJ1f31eKygyd8p9oiY6WeI9zkAEcc1EOoC/2
l5kXc2sLOP5XlvOw2o30ZsgVuanOVkwOj3lHLFAZabxddBjER4NHg682NJRbMCpxVE8OIcj+chf4
vq1qYY96h7EIDgd+auundzYkfP6ZXwqm9JcQTNTmhkPyh2ZVyMCwCWSwfR5Po4ElapRWL+AzNF6r
JkMA1M2e26QCm6vuXsbiitssnhSaQ+nZ4BUCGP3QXtshNiZkDcvbAvrZsjGA8I6pcoUgRhjKYQ71
zdJl6BCjzT4Q6Oq13O/SSgAywEvVzkyFpsKjckI4adk6SVTKJljJ0yiLoz6jADjYG+uJUw17B7p3
1QIWdRa7iWAphkQKzpUIRMby3Ga7TNoqJjm7pYrnPmKcDW1urSF8lmztRlJBv/8ERwbl+/rqcTYz
He/cRn8H+YzOCkRc6TneMQfqsYUYG5nRVMEAVBzjtSCFbbEEPRC+x7TVFPA9aPk0bG816m2QTPjA
XPhBw0I0ClwUZa0w781bAc3JE5mJtnaq3Ib5PXcQ9ZLnBbfbkbiwxGtR+DMfM4aE6/CzwV7LKn+U
JDbTdExbrRS88GOGbsCn6lWbXOL1Dk/Y+/oV/IuyAGbhmqKHHORST/6m2EyAEjOKRLiYOYVRHjyQ
QTNB5iX3P0/Va1KOHoT9HIKtvWbAV9S1yAhZQPbSmUAfuzK+OtuPPNG7xqizdik1Eak29IVDFpaK
0KTY8aWcL6+j56L5NsesiDs23fh33Zju+A2gnMAEaSb5Ow0ECuM7FNJTvQ3Qq2fRse3yl1zx1yOd
1dIUWgfMKtYm7IyxXCMI7UEBTXsH2t+4si54Pfl1/qbZOoFkrXd/SWPGFUXAmmGxXKNuFC4FbDNW
ii86QttR3eRs+8kNmzeSMsgAcw3xA+7UGyZ0PJhLOXgGTu5xk3najMvpHSKmyLEe7sGjxYoHe9Np
UExNYqe8bjKyZag5f/bJyDdCweO6cJWiCQa7PN958ZYXSLuVAjAZDS8Mi72grchpDWE4awLYp5VT
PnUQvSCa1DNsLsCjG79Fajam4sUzC57OYab5Ay4DV3PCyUb8ZFEZoMiI/mFld9zkyYL0nKMEXBxI
OzVEXrTIG3nsTIRsqV99y9Nyh70Sjz1k7D50guIZ+ZI3FNXt8HCsiOxmR95cS3OhaPht1y3pk8+R
ylHyWDtbMa8sPWgpeTEs83889BuugesGMU6UtZ/RMECGfrZLnQLlRhFMcgSJKLOT0zYxot4k/wVk
Icoa2oNM0Y3EPPAain0ZcHJzkQATaI85YBNSJ28/W86ZSOTCxY6+T13Z6ceU9OyOhy/44RHUkPSw
7v9OcchtRdHcYRMhtddiF8Prkxl980JReArZTlHV7ydb/L4Fay5KBZQHyAB733iLUKZ/AOts1sWH
UyzS4+eXY+BnULBPO6O+kquaOvz9OwWxkO+jsjiKh8qXpJRvbKv4uVa31TbVlAMJu1IkN83VOdZN
AifCGf/tED2BJZwF5UmlstovHT8CstBjVqTZUUGbxqRNA3tZEbNekb7+AWfAPFPbm2HNPcMIda7/
SyDPletnKQGS6gA2qlNmZNxZb3wtZfRF+73Lf4X4BzAjiyiLVeVNRw5T9Pkbjl5/dB5YFAYFNSAa
oJTpE1bJWumR0zjzp4JoCfubtGRiiwFce6PSFdHFoPTcvxmYEwlMcR8NlmwNTtIWUuSa4t5AzpcU
nOdPRCldpdIJ+N4VnUgihVJsPJxOzcpMoiI9d/Xp0VVqPCPju4fNC24t0OoWyb04JMuMxqnNEwgU
9Xgem0zt8fb9Bdeq+rWe8WyyK9gIA8A/y84vCLN/dnj/YgKZROx55XA9VUU0R60a0zW0NzgJqlxx
iWZd50EDHz+EKoyRSM2llSilDUFDzWiwY3oN33yNpZm81MfmTyAnZof8nen3UDnrFZ7EmLiUlspw
AKwMJqddkD2xNP05l583iiN/7JxCXZKUW2opsxPABOIFKfQkoNVfGVlcjRCkhUOZhz44VztOeOEy
jCVt7ae6rpaiv7u2TH+5f0Igqqyg5kulZJHD01K1/qcVtexSFI9FlxfnoVPP596XVB4ifYeltkJo
Dmb6c19Y4lT48zKxE8TmNiWfgdOLc4grkvU/xq4m6nIooyYiXwfX1QOruhJaCtvWwZZ2vdRTwIMZ
974RDKrtv4Si/CsEYZTsbFbcX7TC3hIVFomZnZVD/r8sJpEcosm+oL/qGUU8OzCHAf38lYFcn2dX
b2qi0SMNR71C8YKgmQL7kWB7ajf38i0yjMiXXr55JlMOAC4h9jn/0Zf8FDqu42K0YgD7fampNhjo
Bnc6wAjWRmlu0OKqPHt0x4zFo5MHhQH42y3JLsOSvTBOZy3MlBaTGK7yIeSz4NFMx2wHX8B0M+dK
z4BW/r4ycAbJfxekqcPLKf/6oKuwSuG7lce9Ai7GpR6bac4FZ2jXKoGO9FISMX9nmsDIQgLnslaL
VLTztk5ezmSaa/x2DWJsNaNlvVwYyNnMTkueVjSRDPmqfuGGLaNF/tvMvKqCvz2rO0CsfW/w+6bV
O6yDBU2V3EKycLXzeWfrYFN5arkHCeenCrOzlIVw4UNap4PcKRWBYwRmuUxfaKcKbQC1gjtawCq4
9DTgHobYDLjo/2ioD/1M7BaCDoPiVygL3o/MSNLUaiJBO/3C70/TdM4YG6l80TVwUSA18dMdPOSN
v9o3XLrwJ0xQ4m1uJ6l97iRMmjyUfAotYvvlqcsIrOMIPZoWQxT8HCFEOFxLdJClxYtKub8DOJhj
hbzV26eB0ZyqqQ3adqdKZf9OlhxeEWMF5N0+cj7iUr4v7VHYlX+NvBazA8FfArqvFnwJw8+gA94l
xNDNR6WQPj3JN0u5ozKvQT4XOT8xFul6t1ClxvPMEg2ycLUvptDNH+7NqVVlQAfGdNqx4EFSP5bT
ehXBvPZBEEKz2InERsLy9/yJb2UsBJoIAG1cKqtS/nW6mujcf+pF/b9KCFAZHQMRgclbKYS+r/uq
Qw8bmFeKogOJ/sJ7BfYaLwcz3EGCYwGAgtCPZfovdxwTcWpD8m04tX9mZzAZM4algnwJvBAZuR7b
eXyJS6VTRyOQOcWT/OI0O47KmvOkskouhghwsLree08xj9/kCZiw6lEwB5ZpcRBM2MqQBwvAVmz9
52lbsW8fEl7yKhstwQbcRJfNPPyqQdkicpigDSE/AN4C9OSuKkT1Jhb4AngpaBd3N++n5kGNc8O9
+NaPZdWyAMgyLm7yo9bZK/7rdsWY8ftABY+TTKdJyOoxA6CqIFxZ5444KlGhZjKSzTYFREQ99Kqj
MmjF97wR6Vac2gMCN4Nz7MUsD1qijMSzp1m0Am1izPiyn/GOqpomJIxqinAqB9TkXtBwR4fnXGSc
6tKP4Fyb3hTczBP+uP+7+CE2KRh1lOZnRSgV4hqxCmGdU2Nh3wD7T6ywr71IzX9yEVK7FEloHQUV
ZGgvSo8Woz9SoQMPXtk87NVkWf7Z5/6oradHImhFnOC9HEEPcNHKrr2NFFG8y4HuqoPOcXmrnjHO
cZR2lQtRK332Z4Glw3Wp5HeXre000clcuRJK8ngMOPIBAE7bjks9DbaS+fdi07hecVciSHgx2wpQ
aFWLZ5DANt3Zub3I08AYcKii/XgoKqVpz4Q5d4NBSwlOQBQCJvX55mIWaKmbn2IuM3vRP6Es3yGZ
cQ/UKgGIe2zW9WFPCgEPeXX9525fm7fkaRsSJOSOCH+Iryp6EobvQco0EbFPv9jUOzlLcBeyDPZq
tjWDlteP41E7oqJrYcS2TNX8Vewli/LnchrAEkiTVPt8j0aouQOQspGniMzQiRcNAp+zjgd3/sYn
425JiFxcHpgPsCIVp8ZJJ2XRBfa8htYAvN+1/56Dj+Rh5/K9ImTRUHN8PIYPRg/FJC8+1Z9i/DCC
a3u6ssThuIR0jbTXrsvJmxoPZNS7ZFKH6WHqal6327GV/kbttEjywqmY1Q51CLAJMdRfBz5dyFyA
mFgYPxdGWiKNX9ONmWyjW8MELI+BymlpYfULKC7I7zmtqAkiCKtAlQBZHqvzvQ1mwkLbDuYyXLff
ghTT9Ed5jWmbkKdZ+xwdJol6+wk5eNAr9bZJaf0dPPJBelLj60ZTzVSU3/V0vefosT4Vx69x00Zm
byTF79kpEOJtZym7fT4az6VZRc4zDK4uV7krp1XaiT7i57w0kG1XYoRsrOoORgo6rilrPwyKrFCd
9He/P8nOagXSL0jjBdtfzaXI2qDQkKuVN4vU5g3cSV6Az3hqUwrEf2vB807+z3eoOeIi4FWi+5dq
RGyGN6Qr8gNvEtn2swS589+ycoCV5kG6GPxvufO106xFKO0db2yqsV3m8I2ghs8SSvDsHVQb1U2o
vGrNQESHN8D3B50G29NIJ9tNiO0DwZSa+wW2xQf5biU49PjXzUfHPtJGzKA042S/CR5NvPgrxJcL
M4H7w2Gl2JCBmZipclndpGqVSU86pja+kUE1IEabJ70DIVzWFmQtIafIjCTcLlCyNnV+GhCimgEs
6o83OlnXYHsPDT61pr+OLYaRxqChXmd3Z4wFr2WELvV8suNPa931vDZmqbhL1y3xHIMLf0JFD/TA
zzsWBLfBL87TP9BAibIjF6sjdQN4AhdudSM8sd/ORAiHZbNom6fvBjgxh2P2ucxY4hZhY4P8o1Io
OTTJLhgfZL0zEvGd1HG/17xR+HvPrt+s8iEy+XpEyBljT+JeBi+olAPCI5bF4yCjq+tG7dx1HE9q
osGfKMwlYyRJ2Gdh26M3dBGk/Pcw39S2VCWKecX7pNO5alOE8PlxSaXbR6j9F/DNHO45nsCRO2Ao
atS0KJGgKgngjPxNXHOYg59vLQnIZZKQg9CtAf9RiN/X1bnf7NyLm5zB+6AvmI8kdMXyRoqYp0+k
GZ+fO67rFPw/2hG0BzzB3eAxlEpNq0/WNglaMbPsg5GOsEwSA36OAWg+2djsNZOFf+V72bYoqEdz
9wavPFrxCEnVolX/xBaABLSxuxEdXob0Y8xE++topKXzpObJLIUn9aa/TrA0O9ZjTWyTC9//XTWR
u1yNYj36mG/PpGl69H2Id0o/PvRXyk2ECA9HWikLcMNL0poWAXitG7f9D6l1Xy3vBNgbyPlUEF+z
Qam+0V/HIdDTltsRIiR79gW1gFKuT7YgASzr1lvqNWdbkGeKWT/fDOFkWJ4AMSx3YvDTaQ8596RT
17pJX9Jtmu1wvwFCwUTz6PiKiq7DaS80lR0np9bOA/yyyGEy2rsDuxwMdT2f6Yx/O3aHvDCWAz8k
PHQ55983Kwa55rczq4KTb4oHdWXvYUFNnaKFz5U0Yp3kNE4kELB5mBt4zyaCuBDlHGCfu5eC5zjI
t+9rw0oK+Ic6fvw2vSdbRLVt0FksUcwz1IkZBPwi6zPa5oUEnNqSK+jW6V8ZmPMwVi/STQnLEe2e
wlbPMVB1FnPjObAKrOGda/PZcrEFxPmwJsQttW2+KXxdBApWKpeNMaN91WdUsHr1aXaXbRsq8Q/A
Ng4mKdljonmvjz6b5mquPntqJTsZ7nHAcKkXJjQJGK5ox9Q9uc2XSA+6Djv99jhamGecmAEAb32/
KXzbjSwvXexZ9u4k/q2OEET3wocXZbQRc5aroLsWPfKmnpwOKhy7HdAx8uvdxlkTidqKHOukBIbK
bWyIM6qwexQsNOFnhZojSStoDTQDRAC/ygZg4SBozlTFbQxbm43JzwWlEhD7qxYe4Wa8imdl4XPK
35lIbZsD1uDB0j1EKxjE1i8az/9JvWuQvYO5U2zM7ysq2lFNK8qDS31VZ9QrNa8iarvnFtn387o1
U/1ni7HQH0cvN9xfHzTHG0WVE+urKozZcY6p7NJ6luQ0WsoYSp3Bogd4BPiIQKIRdgUkCxsQ3Upk
l1Mdb6Vk/inC//arp6RyXlU6fHZvA7R6VZP4u9tEDj5D12H1uMbJVv73plcVur4shmPUXSjvhecT
c1MohKbhnJLSEBBHswgw9jeHmEd8tCqg5UnT/ElKK4uHhvbbshWGFPLBR1T9iFAJXwqBuH3Mdr7C
QNejdJBt+IYwZqFqXXp3MaiF6mYmHnEpv4dXuR1ApRKJwT/QQqSxz1zw9dpZWQf5BWKdSyn/VrDP
pMIVlPNteGwTZhASEwBt3ZWDGmoiZ5CaamjsYaTzWlaMZS5eQrtvj2GcGihGg15GDLqjE5r7Hp5g
sTLtRgZwKWKTKu1v7TeNAkswEMg+7B2Rg8sxRy1DV5mMJFZ0pUexwIjoxjavmh57irfX/Q3figtt
7H4HguBmxpozw/8GKwInPj6rRMg7QTlyJcZAFbwfk6Xp+0R598Q8iMOMaqpzPXT8pXby756W3kEf
ZPSGUaee/yef10lGOblfWoEwwhWEAAE/OawTE35hAqGh4W1TVfFHvcg/7bLkJkMukVQai0iSbJeX
irCHEci7G2LnuRev9d2ui2sDNCGXjRvlusP5AsxMoyTW+18tvOp3ND7yh2NzNHAi2Zq7JtbA/fi2
P3kiK7ei8ouAutsTblGqL4M0Hc8xP8pj3p+BJCFtmm5PHBuRvsKRJjZZ7FrdZ5PwHdDS5cnCpfs5
5MJ0TsadnMmgJFPqVH435Ez1X0t8Ktpz/pxsvPAW6mi1lh7CBrg0NNpp8xO9qmgA+uYkDquebeup
3HKqit0Y2VYK099hnxB4K9JkXCCOFIKCEQ7No+u36GN5vuCPYvsDQUrLBaSdI983L1v1fGkanSHS
pMROs5U7PtCdSnpyF4LC2MGT+n3JzBy3yFR0SVlIjChV3uFcMcW1smytekXHhzN5+RLyUCR66cje
6vGpWOgNaKLygnkKzStiZO0NQHR4PWCmIWTdvKVxFq4LlJWiiriS9/c/JOy0w3S/DCeL/1qB7U5Y
0F9gsyfM3uAJx37iOdoradQmkEmTrddreZQF66XDR7TY3wp/7HvQS17HdiUSFnL84e0NTMR5ObXP
nDRztOEm97X/ptWZjj8IPKB4iO5NNOvVPHb+/ipLlpGMzwuWfZPY34GLFgt4MpBZzSpXybz8MgcN
RZU5OhzbKErrBxdR2YOTBO3u3YOgx2inFkVIWlJDxhtAsASG9ChNGquZgws7rihIOpJFmpyEMvyf
3dr4e9SSmXtApYD1POnb+TBb7D00pW4y123T/pxqi4TplynmsonejC72deovF8QMP1pFQrpW1ILJ
OTfPXr+Bzu+AlkYRwd+EtIPToZF8m6JFmRzpTblSGPMln+k2DzE7NaQWSvORF1RN1tjs5Cv1Vz9p
lYDPF6x1ginB+cT7F7HG/p6sjWtm1nUa+1wKxqNnBvwO6s7M1vf89r1re5R81TKpUn5cP60UlYeP
ZmFb2kC+k39ybYmckR9C33xnMrF1Iq68gZvwq4d4YuJe9myWyMDtsT8l7DKfc1TFFGBuGdTvA9gW
rvDzS/Q7RYp+8qqV3t+vc7FvphLMyYsp5cxxGV9FBNG0jz4wxBmNLnR4dhBvZIGxqqf6vCZMnqp7
oWECyjbHBob767sEG9UptPwznVesw4LkWFOJNrvayqITCzbLEN15j3HzzYsm3CRnonmPZXxa7nZW
5YkOiikAnoFhXOZIMlgP24m9v7KQcvK4j1MdwE9HLk32ySHcI/IDtZ/v2nUWoFKBL4AcwWmmZe6W
jerKby6bi/zEtk3+kKdorxBI/88iKz6QU9IpY4C/PD+e8g0SyakBG4WpePjLNIyXDgAYW5FvtZZd
Ewta+0s9YvxlBpVgzF67fg8L4/3Q8eZ1hZcT0+ULUiVlB7a4LhfL7Z6zo8szO00/XF7osaOJRWHg
JuVbELGGyCbhi5//xLQYJz5i4l81IIyt3b+cljr22npl+6o1ly2NjYxZzaElfIlZacQm7Gzf/GFm
hPeiu4/PDGyhefjNmRoJZghcBJQQNUy49Y9po1D3ri4NCFTJnmX/bomiiUZ7YZPeHPIPvg1QgDA4
KMriO+02itQijZWF8gaY/ULqsEfzzbPTihHRdm7HIXPWPhfyZmtYX2it/kAlGjTCyrYrwczarPyI
byUN6yI9gzqDwAjmV0gBddMpblVdlupcKMJgXV19HzbrH/iFzgd5ksp9/n0XEzqvJerffTiVuEKU
HWH5qHz9mvvAFIKhUo14Z/ubaPz+ecy/S2Pu2kk+5dYwOOsvbUlaUFdNK5CEMNiFXn4k0SZwCJ1j
H757NLc3qvklgHT6fSE69PtSZyVaTD6miMwli9XJB4qrzeSwi8IlmRtfZUaE4x3IrWwmi6jVZjCu
bi17Et8YtOIiRvp28IlsUv9ef2U+YT0m12xtkmVRakGd7E3pg7B1stDf9PnVpXC8+dInhteLiGAl
r2vdqD44HLI1ZjBKAhJd619UM4fRn3YdUlqCONJ6f/aEgkrW9ONSSmGaIG/yKButnEcE1KY/9kjn
BUaaBW5Mjd+PWxWbKBVI7IJVYolvCAa0umLDrRluu/5MgDYjNDGjh8qPeKPwDgn1qWCzgIKFqlKt
aSeyI42vy497KMw1EWgB1CwyJB8wlRR6RbCMuvFrNKNEmqjzXTyx90KgMXVSIFn8X8rHThQxRJ6e
uUKQx0n60hEbFsuG/ObHhbNC9OANKb95i2xGt+xIFmwO6eYbow6/RPX7/ivdpK/V/I61cbJ5enfu
21Y1JQRpIfVyC2RmZ9rwyiaokKxrnOQ9c/2VBujOdHuR18+WL4XTaA5C3yd0gMI7h7uRnDzc/+zV
mxWV8bXvi9IN08eEKTNGpbNqWXKjsJ0fXge0uYu/uFdka5gpM3+rBYNA3aG1te4/L1/J8s0Jp72O
lZHBKb3+9fAW6fjb7W1eeQqSBof5tBl+lw/lZHi7emiPaURYwEcYd2XsPO7vO4DAKzIhkJ5sxHn0
SM8H4OT4hQItN6xS9DLmTdxfyZIJ9pDoEHuUvxByWNjVxluyLPxfZfTE2o8+Dm1hj3oMxvPugv2O
6Pu+fPF1A+870vBFVa9H8CXRdX/nv6IjGTSu1c6rAwQElriCxw6E81EWtNrPBWkTv0xO6fgyWz2L
rReYyJjKZLlV974FsF5xq1HaeBRtGWeXBhO0IKOy3WF7p9sUmX4Ne+mjFX7KL6Ca83GyTl/WvfXD
KyYNcHW2WJlV4ap9IB7kkTqDlLTvTwJDOMkXz9L8ZD7/0heswcLHh07aORhPAcdeWjzQtqxkI2Hb
Y41TukiiKzpSc1Wj2NCN0p38Z3ben+n5mo9SYxMuRGNUMDo9J144UhiqN0uBGNtIjBv1jCl7vdW2
631WwpGNtuOxXMLnycyKKHyrdtg+al93shojqrFxoTiBSIdu3XhKMkAA7varpJc4M2F5X5s/5qvO
mNlMKmMTrZWtEP+ejtHGBqT7oWR1+Y1RQwrp6MZnr9x9ClqWHz5ssL1Z54GOIF0P/ZtC3e7mAP87
Q34aEP7UXCy9fRttzUjIuAEs6zzMRU5Qj3RW2cKWOLtpx/b8AvHCavVKU7977Nb0gZoisDB4TYMF
XAxAHYzhqrqLOdxSS/ORRkUcIvejrjtFJ55wD7jK4ib6DFuIHFi9OcnNt9lkQHHEHRkTCuoJAamu
zA+5Q+Qmk1uVeD9NX5QXMn/DOCZoD3ZwJoJeEr1yJb9zh9pHcDKLOEsUmhS6qoGp5/IDggR+dpJZ
xhmCVAEf6RAHmLz3G3vv+pUda24C+mPWSqW9JR+82DlmPMdeDuQGrS7qMyQtr5RlXsCDF+r4Mf3v
RBG1CGy2/jEBu//WefWHJUXwq8UZSe8VeIHBcE7iYU+rKUajhV/hVncKWIYzbHtQpcmdBYtz6uo6
Dm9gtwz66yHBgACqRAcKPTLyM+a8GWnId6W4NdJshNz+3SDASun0IpNpQ7Ek3G0iocGw6mND1P+U
oSu5pQ69g0FyimapttpqKc7I02JHrERIDAgsKks/az/iG6jdu7WpxPWihFyh7hwdlCiQlvaUcyJ+
QTOMMEkksOI3JcksnvYV6ntlL3S805jZZykg0hUfZWFrWpEsFjm43iXwzSrAG/9fpiiGfPnwalD7
5APMDKnX44X4EcuV8WcxQtIqoVk/oXeCPxqrbHIKJEz7io5hDoow57ome73Ify+knXEMFCKJpCiq
zOGCPI2gMosj639NuDfgiSgGgiqLMXe0wjLeSyg9dA5KOLfr1WJOneMaypHFizQ82azbAjbniwYg
Ro1yz9Q83ymx25vrreMfGe3oioqlaKlM2qK6LB/jtvGDgFYaiU1iPUlGK3RZ7R89OdC62/f9ebsT
PRM4gJCnqhxXy2eC5oVF8Dk7PaHWtDUL2X3Tk/vzIUMOgis8ZI3rAK/gzW3qZYhrriUsNIqCyPvt
F8nzu/bQe5+0sGUFG6ZQfJUkMLM1g0KrXWq7rOS4wDYuHxW9CzgvboWuzmmitbi+Sbu8b10aN8QG
iI0PCWoBSVudHboOwSjLbITwEUsWYAK95WBCI/LyArvJ7/ZxJQ8ls6JpfCnNQIkEakHQ8H81Cy7T
yfIJGpGPLny+eVkuf2AdgTa+zBefilnUVD3ZmZ0n4UewigBuWOQUbml3VWMbfq5deOV98uSp359A
dl25Tq73TfBnZjFd+MqtH03wKWzIwD0q1oAO3sKDMvf85LEfSucSTVjAvQF0OfTjj41kGuj//xtD
VN+Btx7XYCJqTG+h31ygJEuGlhsUAiG0wMjic5vN8xGQrUSkFEzbp9X2fs2ZToYEjAJTFzejjhoH
3WZrWSvmX5q6wO9GgpKrQvxPvXkeJXiySyixKI+55CyJSvZhXR4iQ9xCfB+fO2LHZA+90J1wj70n
IXskdwy6SvRBd/GA0bxcNCATTjAF+vSKtswA7ylWp9ZMIBQ5kcq6jx36ySlOpCf2dyP972GNKIWb
pS8yXpqsl21d0ZooJ+jnyMC486vbRI1isvezL6GtrNmr62SdCWPY8UWlLSIMUeCYzF+J5t0RHsR6
fleApEFgyww/5OMCNi3G7YjTXs40+9R/Dd07n+MegXCJfutTP6ul8aVCzJ7NAtKftwKVtiE+fBNl
y6TD5Jj52Rl+brOpmIiHPLvOnXcDjpFUl/VubuqxJFYLNhbg0mRddWTzHq0s+Du9610qvQTznSY6
Q9bHJOsbakNHpr5rK0SeTxQ52X0UkOpgxHHSIivZKnoXZ0GUhdMunmMrNIZBx3KkBbNesNKQ+E10
dZN6welfQl0P+joruAQyd5pFCYAFs2gWDKGBHRlYTtqK6pxb/En7AaEn6T4isHFjxGNzyqB/sz5C
JvXX5yEPabGeyC16ia3iYmt9j4qQyAizhDt1dxL2iDZBg/hLTYlb9ztLqfkTtpt4F/GoE59xGaQN
JcMVyYwCExtbGMdUAl99qX+DzmMLbG/8+t1LffpdfpqKuPBdIxyNau3ZIt3EJuSAPkfxS4ZfUdVi
SxzqnHv3odHpdcZSkiyq9+Urbr4ei7SwOJ48SWtsSCET8YCChauAlPSW25bMadroPZwezT7fLvax
1LV/+fU61rWGa9daSxl/wk1CZxgted716zvTnAarmS9kgcplAHR2ufVU1vzVw1MUbEQtDfABh7Zc
iizTj4JDoDTWiV/eHu895y0YWDF4Ujav5hD4tqNI9x8F3gPQs2GNRf8J7LU4rFwFPhkUX3REVaww
Mum6WW4w4LSMMui/tG1QRjJNfSUXcz/409n3+nTDQY1w8qcNRve9k7WKCtSXh20tlYLDLK9FsV0M
joTVEcSgPzvztds9fndlWQ/F+968B0HtsqupwQu3uf463q4MddvI2ty8VH+1haiqgxRl71QS99oV
d3le1F6ltrv14vKicofeD16gTdoZaFYXMB+O/SSAl7lcUAPQQwhiwCmC8iaZ4QxF97RTZW1dR3Yz
RjpqupXUtgXlFGybUgm5iJAg7tBiJDZiOE2JjtutIiXlSDQ72OY8cK440SAlAW1izrvaHT9+evbY
4VSU/zlrXACfLValZibOqM3xkRqkSdadLipiT7M1C87fr7PzOta5g4nTi9M8v4LM2DPxDvG9CmHT
CVkW7XwxB8WpGt66Itu8F8OkkfMObfGcem+xyoSYwFN2Zjh6KY43v0CDAb8EfLFQLOqiYg4F6DRW
x9lJsNcgYhnszApqsjg0tC9yF6qez4ksPQdj3nDn3COIneEq5P8BJXXjyGWVCCocGZKvtzuzm2FV
6ml5IgPAlLi/DsQJ7iTMrcpjRbqHyZ68d4w+yRSjWFQfhVcXspv2XWS4bzbDs87jGu17UyQtBhH3
8aLurLUsvCiIGzoQAFHN3UaSa2UiLD6bIa8CBJhjYfnyjYhZ2E5lqRfAFUiPWqp5pgC6DCB0Cxum
nm5LCyqMGtmkW8GcH3LecCCkab4obxkeOFLKGFL2yFk6XcKl40od9g7saDRz92InFPHI/GVvDdLX
IZSzqba1MIWKnn0qpbcwOxwsaBScN0az9D1suXczyMxgW0L2CBHvM0Lb+SDJFKWYEwogghgGHr+S
dkzLKcWpP6Qq0Zy9hCz8MYtJzFdp+h4gC1nDlIxDWVZ9MbwvNcBfxsvW0onZiUau7/6kYZblzR6n
orySoAdXBPEa3DodKsAtj4buYY+eiFydjxoRe8aLJ1g8942l/K1f2FE+S3rY0/vgZsGnU1PoT+2V
XzlkbMITWB7I+HmiRaB/wLItiZzGzUyTKaJL87rg2ZXK9gWkc2/XIsLyC41BADTs0tcOAHJxc5a3
9KGB5nN0JN+8r5gtvFt6TJtELVgYjIaNE2MLymAxIalM4nPELROBWdY+uLy+sVIc+id8GoPK12d4
976S+r26fpPVTeHQGrK5jXgwRipWNzFnNN6mDXMy5igZ0ina9bTAH1tg0g84b7NCCgoGgwkwecLp
HnawgvgGJhw3MBdh5mctwmoSK4v21zscHnQEdzS8MB34idjbHGA5wOtM0vIb8+2JpKiMdpR6KrRQ
TqSn3YLIHTGuJlvTU++5uIXpLQHUuTwcR3MqqLRTh7Mk3eEppPuz7IuYNLgGnV1dfI50TTINCbh2
RS1KJNxTu3JhTJhIUMBog8no0sEb5Vx2rKwTch+OWGEl03hsp2GH1JUIHvQBAJ+u+SE109IpIbw/
yKV5EEnMwVwo48GXKvKsfcR+xE6yr2aGMJtL959QyOedfwcgi6GHCWD7L1ibogpAQP62GwVGqnrZ
FjWl3mZg/PteYx3fKNGo06vY/lnipdlA/s3H8k7/EaRORV3i0fikY2voaIzJA/JflZzs86xX6Uaf
gOVpFVI9Iu+ly4qRimf0BjVYyNxNEUck+aWe60K8Rtiubey6ZsnSkuVjSiFcPOogSrvhKJLInvxY
jweroMrEBIty7vIN1kGNPtQblKa7RjVU2kq8V9ace4/dwrr8O5Ey7kR7ARfq09291baruaGEdiwF
ghAA5qF8smwalyUFJ6yqxgVPkY9DediTXXZ2TrWmN+cIv27o1KmqSjijuy74TGMusKL8AXVpFLgR
d4q9cz49rwqGTnu5Wmawdn/xLzSTw18Iuq+Z+ABsywJYACivwO21e1ZorsyeKuBUbIgGTcudvtMC
E1xBMqcQW9h50YIrbN5djYjsqQi2kJ8Ne1lQW055U2oJ9/C5ks0NAkBnv1nAA1NXT/z9vHw8MmWw
X1yFm9+1mcpzsHRob3lfNUSJd25XRfBf8PVcp0VwUVSiF8WJPd3SnfL8r8TPiIxIanJJHM82PFLG
46Fu5eTWHfUirufzyU82BUJT16dbE5TeMiTqSuXtcIMVnt9cwmmOb8cvdUC8oMyu3xjk8uQohtg/
Zb24m5IA6aa3YGbdUJkU2z4zzxv1+acE2yqzGRiZQlYMueulE1sXJLUFVbHdFWg/pYGIBHnHH09s
oM0pOQKtWkLmHFWpKteoFHlcaAx39/cwsTkeOyNz/eBEuHtjqo1+aipeCgKniJIMvWIEpIIIgSTe
zoOvgoQ0UXoGWy7wqolsYgf48Q+472gFcaw7/ArXCXke+fGCImh1td3tah/IMfNngVFV1h69MwDM
88tVAN5Ic9SPTLN2Lbab+oBCZKlybu7fjNJFn6nXcW9O/kxfQVwwYPYORVcZTMTPIKWGlL5ZA5tB
vXsB30PqvGwlO0nuaoB42i1YCLFFltGuZsE3TUPVrse3VDWB3llr40K95wkWsdBkXAQqKkDeNzf/
7Rxxl5KlnTxsJQRhmu3+Bmo1sMo0QzYKvuZnHF078FdVQPmq/xSm0wEUWo5paHuuOsPdaVmgjD0e
gVj9QZMGRGkWQKr8e6A//0Av2NjKgIQ8GjfQk84A17SCT9CJOHFm4oe6tGo1U3ZUdzEijdR1QXII
b46H8yI6KNOrWagWC0zdNUcoZk/8sIo8xEaMEwC7zfExvu1JSzpypmYqVHeuqtP9yio4jQoYSRlH
RHfcddE//ujq/kWj+G28b+6OC4+vJKm1bW0JReSPmgyzesTx2R2yz+dUIFgVywsxz0PWZ7WXEZjr
+8SKmwVfI75pVSbPiGjNJF2qDOimS4F1gf0xdLm7JdNwiV/thlATCP3tTJMBnY+Pa+pA95hoRyEa
Y5MpNwLpqBXFMpdkSrlxGRARvOwfhYx/PIn1mpP/8aEtkqZZCH7rG8duJv0pio1s/HIELdWfeP1i
scTHKBSuKSOMX6Lq8cdf/p2fZscoQkoEJObpUUfl1q5b+xuct7OSmwz2m8m6KdEdVCxGuhyTV3YV
sgZbrQpzyOLpHAchxYJynYUTT5l/iAAIwdxcdr2qWAHmZumzn/6p32plJM4hn2baEh2Ov7nMb8GC
X7qgPA8RB+1isE+DyWyvhV/gWNcjl08C0Ki057D7ku/LEwYUHDg+svKvlY4s8QV6Ey9ZkwIs7R2D
hJxeigxwBt36CdiXUQqKUL/hrVFmKgyVcormMhWCHcPIHWFaJoOoYw/ljQI1wGyPI/GdQIEnITQc
w7+69XioFa7IWwogrU/+pd80GiEzPOBfi3Nns4KocxTTHH2WkdGvtMf5gbXMPLcmJ/gg0tEsBtUk
wwqpmlEp7DTSqZaPOopDPY/d7fceoa0mZWiBg6sYF3C6Rzfx/uYi0sY6U9MP1Xpz3W6j8PyHfJcQ
XaVK1zh+G+Wbu/SdIDgSCHFYzJQaSHJys6YMjr4JJ0EqNWWIsg4pDd1t7FkYkW5nXRpbVCOieJns
4qK/SHd5sZC1DM9i/QmO+wTU+oTM2qpeJkH3xDphz6nmDYsT/+h0PXajis6xnJ2Rvun58/E1MSuC
p8toVhr5YPDOwtE7LNVL04FFreWDYrOVzgXgknKi/G+ykyAmXBrgh7BvubuRxcW42NVHP/AFzz2H
erP9ps2DUE5HkAGw4cQfYr8PvRa6nBHkUTafAR2tYgmtN//QSK97kxeJ8C5m9Amrh7v7ciJhd+gD
INPX2hiHKBkECOsFiIv5PXkPRiiHT45hw3A+nQzYbz1eumfb2SL7MQYIXoA9QpAyxTxyruYhE7f8
hCqWWBtdyaVfVKkFHBcZtPHnj0LR2b5E7GM2FDOqI6OudKsGeQGRWejgSH9Oa0Ek5pF9cAe5wu/5
fX4P2zt+KM0zjJ3m28YcX5M2nqPaYAAtMxq+0Hv3R/eibAu/JM66r/iRSK44h2WZrE6GBvEcynD/
TXO1mxErYxjaJ/EXFRp/DEixFQztOWHGek/09RFgWUEEnPicZD2uUmKGQDXSHpz1ehPkKuaRWF05
ZBFxNuJTlKwmmGyaofF0ynYV6c6N/DBFwYyH4fEjJEU9+h/6sDhaqLpl/IAjK/Em4WK8D9d9ZH/z
dr4orY20d6rHFcgkB7uRBhfdvQbESAkG6s0HnnLBtYSonm9CB/uHp0EctbAHTd7fvWnlOrlyQq/o
+7v+9skM/xZHT5eeV9mGULvEf8g1YXcVtUke7QPoFyUd9jpw+dE9b5SYB+69vluQyl158FUuw6SV
Slu/2SJNcwTI2MncsBpAyUVAxqXEHOdrlSa95pHT53lmYALg8jwsoeDhvju+CZrV1o9zpp8X8p5B
4J1vqBW8CowZzi2fHYDUp0CXD/w4TzqL+mCE0KWQwOVd2opddZ8IUCSJsyy7DN6QTUEfA0R+1WJd
98ko0A828brmVkEwgxrTYmTHtuWqj7N/Iy/B2hx40xNKYOhEW2Ro/MRj7lzSPed7siH9+pAbDYq+
GCE8OVakY+EGkyB/ybF38JVxY9OlXU08YVlKgh46JnfvK6GhFhA9PkIGYXXQ/eUt+TdegcSJ1PCj
noZO3gqrFCSKva09i8/ygDIhD2I9HKlz8mbL4G8Ni9LV8eLktaCzXKnn2ANIKBLfh07b3SER4jue
aOwHf6MENbBSU3rh8JocQZrEs+ERHLdzqcQjmZS+sh0Vs6wqQhTvRL0k0wpr1vkgk9HMWJePQoUK
payDqweO6xEKss4Ro6KXZNC36+h14q2qn+VQSSXCj7zrwf1OwVweC+HM/E1lMr1seNmVXeYvmoIc
1w2GYkOL3YWmX3u/Mj+Sn0XhFOTSLLebmdhPh7YxjWMFMFU38Ys6ozX6d2on1LTgmHNS93ryy+EV
/db+FhmLwDB+38SVgu0sCpLlvd0Ch7+LJX3+LblNhTrIY2JEfnpwB3qaTova9mOYvr36v3PSx0nK
7Yotkb06IZC2vnWBWLLURAsNhOuWMOmMKlXEbwKx9j6qOQQj2MwPu5JKL9C2qeCoNuNv38wIwn81
5tmazZVdRV5T04kqrnd0p28Pwu4kQDOFilALd7haKeDKM4sYpgQNqwhXhktSIvhwYlgxcrvW3j41
w3Xnq2NSiyBIMAKyGCZZTESAL+JahzlLJOMRti3S/DAP8AxI2AgK+3WTgjHICYzb310B2P7gu4iW
IDAF4mr9K0Mvrn8xDEAYB0pKiAKPcnVbbREXixAqKbyRigyEhpmoYP7TALdaeuv0nhV28Wvmng6i
65dz0EnsZPiQQE52MeTwDoItHmwtrFY/AQ7nNqZB4RPXHotNuRrm7YnGnvg8wk3MOOrYVeoirVuj
hDsNs4YFHVYvWtqZKdt/cG/wnpLbNgIRxCXHg2fr/qOJOziIHISGfVDJp08a7rv7hBEKni3bVqMy
vgBgTt7AI9IYQqxN6o3Cd7FikidO7EiHsg5nIow+1q4r2u95Yd6eY/EwxnSBtVnSAX3tM8gxlbxZ
+lzwf6jJhXPH3oHrmfwnblN44LgDOA9wwxWzF52b84fvEyJ2Rh5b92Uk9EYpUsw5nzbK+QkeiE6C
nmZfdhoJQRJlg0ALFTiF6GSrri6ZHmj7CwLYlRLsqqzfHPRpfmJ3ZH/I78Snvd8TVyKdNxHw2wNX
Kod2yoLMFIlcelsXzq5w4+OceV3mPNX/E6xbulS5rD+DWY9m/ShAWm0oJfTHN2uqKBhsPoPl+ruC
N8dXhJMen5u2MbTb9f+FhPph7FY8OUz+XGWtliIefwx0JC0IGP9Wt3Lkaylpmts03oKab935X7/6
pH17YhNm926KBiZE+Vr8FJBxCmfrlBB33yFAfDgiGrTxWtVAdH+PuQaGitQaC+Y/30uoWEpwEUbG
/fDaCbrS7lH4kZXVA4fcDeKCFd/XAqQVnRRHDk881naY5V/lzhUhUdyJhXlLHAbRwS+uo7fzz6MP
pfUJMztV/R3VNQS9cUmNcTVET+ab2YUOUgkgBWKYtOspwvchLuk0BmRgbpYGq2FN1e83Mnstfz/L
EoMiWyh6oAukvMVGaMm6MFMekHRDYxBC4SX0gbeGYpf0kceVhZiRyPoI9LDipbKsyjPdIZFRY1rM
mBT16tHrUu9iMa8LidTzs5/LNf9Z2kZoLnR3g3dmjQEipihVmChHcp645pl2FFJMZq0gyEy+foxd
KwG8rXcGwo0a4nRjC+zzj6aDRjp4J+2KHBNbM39i4ui3eR61l3l/zU8NfKlw9Jedqv0+FhsjlqXx
QwFnvi/+WUxw36eVIljn7XCqON41xEeG5GMVGCz42e7JXws64lj9iWqLV51rEck0gP4O2OpYYBqz
wikxnv3L8myFO6yvgLVw3PYac95QrOjzu/lSaPlfzGigtmEn6sa54CAIOWRhyV4gqPi/kgA7Zi9e
HlNTgpBDAdfcws8VaBrcdahgkSanryjG9sbOBqEdqjOGrqJqjzDSNipkvACGMFpHybHBfTIa+qzD
NZZlmeU/pB9mryPqIaZBsr4+RwmvPPzXC2qybM3hhSYcH4uk9X1Y5luXM1R6v6LffxIa9w+UYk/5
pG2nEvxQ4mfF98E+tLLlwimsLNXTT6h43MChAq4VNYxnYc9Sbdq7Hn8NGCpU2S/zGHMM5skHXieL
1qS69143yefoGifHtevW4zpyQoSoFr4Xho5ANWqFf8/7QdGI9DHXyoWAaiPGmaM1DxesVFHDkwBs
ucTg6T7G51RHUbQpgKkpE1XtfvJLeFhZwvRP82pANcXryfaejz665ZpdyP0HGt77Ni901TyFt6oV
VPtoOImkB/sCtP+h+KCPyI19HYv2hRIKlo56sL+JtbpzXMYSbWxgEcHWGQEAM97Xjx5EnUM2EeBn
48lLDl88D3S1MfophLXID7DNH+IXxGiqG9qiAb9GovBpI14fMWXQvuHmX4Yd9011uYeFu28TKCQD
VlzBZRImgkCgs6vv37cxXUTPizc3TmGF5BShNFFVj5efCHgtl4XHD/f6c+aWEYoMvMg8ygL7rWM+
X9gJ3+d0B8lqdQVAgYUcDcd5DNzepBmuSD0WOelC7n2vnw6/sVIhokJPzqMGLr/hA47WFFOKNWCk
A+KjJ0+ofPDO/Imgw95Umh3iN/93GOrN79QrYgAFo1g7iSFW6ZbiWbH0u5NJj0Zl6IiCmBVAJy6k
qvjJz4RT474UKKe5ZS9VmFhvrlYGcLydUYVh56wCUJZAOt1k2yF9wcNoZ36YkQXk1JRyh/y6ZX58
iGtDD6s87kpaKhxDV41qjlFPSFv0iMJT4psJ6DJ/BVNdJMw+VBuQPeUy266elOYzj0zf5kG9nJhU
PXjbduCeGVMkAfQtYz3jvLi8f0oF2dvO/WtsnmWPUuWuihGRIqzhNoKl3N4a3r7HZy8zE6bpFy8C
GAhNO1I8S8Y9+jj6nEPQxeZ/Hdvy/2PaSXnLjG4i8GiJ1gz396qJo/y0CUj0Hld7R/PUtjXY2MlK
ySk9vKQHCKfVecrCdIzHvm3Hp5L9Mb/znj3yLKThppaeQ4ZouJdAnh1W1M/DVaMkF+pbZKdWxeeb
R2p4FVysyDyPE2HwLDkZ0JRc/y2lvYFmJSWu/bX4qFwemaPNpSFlGnwjFbmLIxrmqtDshPFlHsss
epnjEJe1GdHSu3uYBwCPTbJ0i7Vc8yzRctu5CuDsW2WAg6/KNc01Q4aK2Aa7CCQPr/GETvDMHP4V
3c48G88ptAS6uYqdR1d52PhkQo/y/FKNMheQhB9TzvC6OuNTRbpNmTiyNDHA/vPvamErLc8raHj0
3ND3HlGuAZ8k5TNc6+fq1RVwkXMZcBzAQh9lYwXNPY0UogqF1/MNoNFvfiSnwQQiOsR6AXxX+/aN
lzZFn37EmKmyOftfm6VscC6ZqU6ceI73ZL9IUEK2aU1azdn23iQ9fDF3mFtTWM3kcP5K/+j17dVi
giK7aHlqaDRCBUdNFjW+srOvajRXpg4YfP3J5zbgZVeikRwKyDkCbKpu/+sLFbwRlTMtvZLBn3hz
feOL0CV6WnZpEgEhUsA09T9nFDRgF7Z4IkbDrn9uIdeMpXK+ffcsYnLPJs37jodSDXrOGDFd1ufG
lyBWZqZU/bhu6LRKVY33HRYOvHBOPnLk59rJ/doB6JcAUP6Z6pVVGJJW8M6Kh5H5ouKU9MOQ/JQk
AbqTfipYi+boaxhDV9hHYamqEM1p21X57LY8DTyN31quf25xph3RGq2OsO86SUuE5sz0qu4aMOqE
em37L3gOwGYa2itQD2gfavZpmpbl1Zkj7+PdQOa+AbR+I+xdvW/wA32TUaZbvRicjWADRS2C4CCe
7mx2e/KFHYQA/fRx49i79ra8EOkKvWWMl9HE93wyDA0PnB7RF4C7+auaaoFbSCtnS2W0GZ3gxC2V
vo1cDq6pwu4Vj3uwvUw3jinMpBtdXJI4Z5Sqkr8uPvitYi9ArSPkuB9CVktEryoEnZCnublsjphN
63q/31T7f5c3RV2GIfnPNc2QTQpcnZkBCUJ78IXodqd9lLfsW6XOWlmrFFjskKbtnaLxGyB03CLA
ubw4ziGeZ1SqViSUo1OLCbXnqheZ3C1Aiomta2jffx8xQ69p/v8BY7d2kVeTVE15BYDNi0FnqMbq
cMOwmxqwcnVm6tnY2SH4FsokR0QnVaPJHtCdpoUwe+76hl8xiqsJ1eH4b70EJ5WbALDOkY5pnNSQ
PzG7ss1xgLeajf6tQr/F0y/9XQhA8VLNNKZVypzbG0cHaRprofJZLoTGnIuduF0Q2n3Vmha8Qxa8
dNsaMT0xikQvBjM9TwRePZ0ZKSTbh+VcFIywuBh+xZtCnQ2yVuYPLhL0UnjbP6dCidx0Ow9eeyle
05K7fPPaHg8ySDj7RR36xpVfUz/9Oq6ZzAO+uYetgLa1NotOjhIxPP/HSPEFjdBBzdxFyRKPrr+u
G/OyXasU2CwPYYVa1lAt2U5kaZILqJN+4sYfU/IEaJGFL/l5pwiY7/HUPfmgoDdMaOkKqIzj3iPM
YCzA0pSg51bkD4eEXAyGsb5AH+yBBLrLX8vP13FaCI3RIgONoS1HvtNzPA7QXhcQsyaQvzguMv8r
Oo6nwtM7XBW4oombqctcuXswnJJNqyB5gwot+wS+spuGSSfRSXEIEiWRAEJdRs5Y/AsgzGoHMnYL
98MES0Am6CtWNw8UZGq0H4DKXKMydJsyl2X13JdxQfe/8/gjLnuUc3ghLYuF9307hzvK6ybZpxdt
Yp3jWfniJkJClH7zIPPUJVVBQ2g2vzrjYAFZv/B9bZJ17J4nzAwuuN2+KDzEMsKTofZsDH9u3vFT
G0wxNzpJrAOrTM0nF3PduHeG/RqJ5TI9Ggq/COaPxHVMYPZVEoymFee49k6aM5MCKaxC2adytlHm
j9H6lGGcO/5nJuWNXG72zPYc1iC6YUPQ/JQTjr+e+TV2F4+wnEOiOC5ySmqP07tTlX0+Nh3EkfXj
9isYTGd87MH/d86UsNjtML5dnXygBCLLo+51WbbeIBvzrP9sCJtM4cBoGh1+7E8/FPKcG5PsERlQ
27VqUj/v3z77gwSWXxdMheZl8N0jc+dNL9G8KF1aPWiguMfF9ekwolvL9ySz8F4OdmfIv1QOFM6R
0Mu3EYLTlQ0E18aRKBTQssKYVtU4syPYjUrj4tNR2T+HzpbVaCrlKIfvb9Nx2cUmPnI22poSFVrR
Nw/orHHtOsDKlumotXB66cl2l2iN4n+QBKtSC01d5U45ycLo6b76dRpIzY0QRFvRv0I6rR22M/7a
jjio4WJxoaybC+1mkGHOzH00+myysADsLTwG0jfqdmTVqWeYeNWhyGFVHgvZSXHQskaqsplzDj5D
YhzW1d+0tC3oHB59G3Mb5+UZ8a7D5T08vQpeH9OELWqRidv88vHiLlrq0fg4qAXSJAY/8gOYlCFu
PkDKooQ+Kmdhh462d4DOfMqkazUTP12em/53QlLYErbbW48LyivJo1flLCPf2xmap1sAg+q38gcI
kUYvQz1wr9j9GDFn7sq5x6OIZbHDNyo/3Cu+LpJyVOHihVd9tc02XU+C/ZiMDB4w07hvKdxayIME
Ow4ZN0yWumqmfnE89m9yA+YuS04OTejtUVn/ifGB6tfNt+fMWeYySNQaDtKvwNFbLCyKYnDaClvY
O5FqHEnGv2S0WoZ1KOhRgXccDWl0CqP5yjGF9rUtve8ChKRr3mjXHf0AAKpatOdJeFiGVDL7ed1U
UPSI+iBgDnYxrMoiOmzy1NejCtmGlQW/XIJU06zrr7oTb+Ji2CBs3iic/LfRJ4qJoyJUuIfF5f68
dH5Pow1qsd6LW+IE3ujPZZ+zQj+NlfVt460zoiCmKirTbH94XlTiiXk97oIqf/KWEl/BwQ9f48rN
cjkoxnShA8yxdIsSikmCNxWGZ9YHapJA8NaFZHkK9CCImZfHeY3e8dPHBuUdnERLlD77ihpI3dZI
9ePrSyOn+pn9gsr86LiDWFuFptELc7Kh3NQ7IMs5fTy1GN0XTh6TBseQE1CwWt4fr07KIrELaeYJ
gMzTnxKerhbNny18YoWmwdT0fYjphHPhyZ6eE0s8Ah1zOELpWjbrlmXKVm0jBfk6WM0cMQ31+rhl
64uaGw2XcZXcgkberhXDff68f2XJWF2uwXRPGIlBtZd49JzNQKufUbP3tPBEuHTXCPys4bCddLNx
Bfca3w+TrzgOC9gKiCAN16mPijBvfmZCnrGAraGKVVptqtSykTC2voLCypN2Y1f3edOr58fHlQyQ
Ji7uxqxcrwyl3+MIDG+XNBY90EO11NqLGBAGwTGu4Ac9J+/I+xiC0fLkr91cv2IBG4psI0n2+54n
dJIjaP3y1+SsiuScr/KuAXyW/vlmufOftexXFnjxZweuDonvRsQ/YrZJK6iDxNo7w8DbMO/Ix43W
uCp1yodoJtbIloXWH0kHiJWH3u7YB4kF4jhIXZxe7gyTA1GNaGm+pejOazIP2fW8gQYZIiCdommH
l3BysmpYgp0Hsi7unCIRblGlsIcjVt3hgv7wuUzfIxbyeK+Ivx0hPSrOFLa18TjJMSFxvPjpUYpD
PhbViXRb77piYv1rUItw00zxzVd4DganbtPTzJnsZpFAMc8KtrXabJn1WI0U8LChcEnzF+5anPHi
kKeQwxN72tGYKWtCABq0TBLuP5y3ig4VztfdCgZZ
`protect end_protected

