`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FqqmXG2bmkDfgLFyqWtwC7ABQJhdhSxfeu66JE1xWCDyDQ3Immm11P2o4bfbxkWqoOyvvCVIKgLf
5b6bTG39YBsYwYdhkSLmdTPfNlvliF+m+KFGDhI4qCvGDSuSK3kO5WGn/ay7d5fbjWYotyLT6Xoa
i0ifkNLl0xc+IU01Nt1/MRCZVwRRPTFevGnZnHn35SVdznZH7S7b6nZ9nIDybHope/r6G7wn1M+R
z9dAL2r3kA2if4gTW6rpLJVqWQ8S11nAycRifDzkLWf4fn1M7ZnvcgGVynY5B94euhZDhSvalYPG
028pjIcXdfjr3qkC1YjxYb6YELimrhLDjZnH2Q==
`protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`protect key_block
NRd+nk1olTHcHRokoklVVoZFmI0U/sOcHu1qs1uCioJtRwLOGlEHPY37E8MYV2zCC+vLsmqJ4xGU
TgHxL2YRXqVo1b1A19OcujnWAO+R3i3LoowO1IrVGLIkwjy9C3mjPymAJbzGcSWaDJscPOVX+/tE
COioFK7Hsv9RG0cG1Cw779YfzzBlZfzmXUVogsoL9G8zn83tN/03V2WIgnCJGc0vF1O6ssFT3aHy
zhjUthVBBiDVWXnRBGfYtmsLwoqomKtvcgKNjchpputq3GXI8D5ZQKMlb6xcENmkdT23uo0cPthb
Tyx5ugQmWyl7L9Z6CNAXRQNdaBo44Z4KZ0CtjwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AQrfXTtytzZJe6QzMWyQ+6rn8yNn84eM1jSJTC8gW+LuoQBONwrUgmnasAZ6xWf2ZxqYJDxYTEo8
gAUt+Grs1g==
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gqEV9GAZEOcG1xfqfR3iZKlCZ3dSDOSPVeFpuBLH1Ns9ScWoAc7vjii7bCVb+iNTXlNSNH9+A+hN
s4KomGS3wWS49KmZEFGUWfWpknhcUgcLDQdkxa4W97Va5GymPFrJf1DodZ7HOoeW/5enm5UVX9oa
wNAC9Q6XZRFPW75XBzCaM1mXJmJnoLroLPK1UtMVkqqtP/1mNXSwAjTkhWlZGT9wQyTGVAzkfdAJ
c/qY4YS9mi6TJGp7bntvEEkSRY/tNOYWqWCPB7/L7q7HOJhagGTD71Q0yvgJKyjcofaMAcEtbxdT
gpYROPj02zQhH6/cyirn6eDKffU2M7+7O2km5Q==
`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZVB9c9OUDVHUgT44DKMnslV1oXwZTtVFjOWqgX0NuN3TGYHBn7nR3U0dYD4S5SN9KtIy5kCboWDr
Lff75vjbFEi5xXwiA6wN9HNtzqkKC7VSDmUKJBp1JIvuXumnZsSJdC8PF1h+yYWcyIp3NtUiuTBJ
6wYeLF3vmB5MeuRo8WtocTlPe4lLwWthu3ppxMV19U9NVWETEO6Ivq3kIxnsRP4s4Ulxuo2HRAOy
6Y86Wa/fAvUvZ8ALvcaFUoRJUldPd34qQG49YL5FAP24fE+Eyf5oyNYNsisNKi/gVyrfNg+HC06z
jpcOQkIEH01Kh/yfxYkqLijWzuHFMWIdTzjxQQ==
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bQRPd7ECXKNhsSUTH9whu+9+6Bw2XWT9ag7mU4kaItvsqZ6jrS3APKMNMmrOXIg+wHJlsQAJrzHJ
dAQPPlWKZl7pIuqXtw3Vk5hlPT5a/6XZqV7VREbRG+z9rRZbQLU8xPFMeYBAChqbB0ZnH0JUbeFT
GvvdGVasqsBxHBjB1+Y=
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O6BIBU5A1i8Kfcpj+cf2yOu1l2ow/ej5AOpagSMW81y3zaIqRgJFnqfBncA7koWQ2YTNRMKEOtHg
bxrDLt6/zyVc/5lPD4ozwxRdxtvnkABNG8e6wZTCMR11NZHERwe+aWx8N6qaLwrB24TgORGZ2DDt
GHtOF9Bl0nCRdW9ZcrpUpi2ZJLG1hay0HWqga8ifs9JUGfeyGszwQUjWHGwLG8QYKTxAX4oQui5V
IRz+CBxi7BjIAlVuEzzaLgKiGVAb2blTRPJzBCI2nPx4PNegKoi+GGEYqgtJZ0lgplPaJE0aaV/8
3KUmkxEhqFR2M0o4+3NcVmO5gWht+EwZh9cGNA==
`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sHbv/24hB7qo55hPFj6kwFTL+oGf1Lw+M0Er6nbK/Rfwc+1bdK60+l4ZLNYQYUjc09CxVlgjEm1k
bHCHAO/YmWFYh1eg/wkGBB/WMKhD//nOHDwGRwxBtkWVBQSW+31rdZoVZqAlam7fwTPpqjZ5h1ES
4USVVx+iigFHouVUIPwWpjQwq37B8/GPzO3NfAMFV4bY+J9+ydFodRbNWe6BX5enTKJhhkJRgY8w
u4nXioU+NUPKR3K+N7AA2otqE66D0UQsQVVIfUvonveSVNoZVhnJ/tk2R9MKfzloU9cDcZeMVr/0
lGSc8ZDaPND6oBorbTikOeHVaaENZvK8wUeMHQ==
`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
g6ni1aj1TrjWZyBlXkgkop04e2TlY6gxA1XDE2PsuzAn2EJmHQ2Mip3rou+FmFlvvVvOTzg9DHeZ
M7a2+ox+otBLJooTRgB1HcYQAN5XiSqXJtHXE2EUUZyqYJyqUivvpLM0Doh4b8efmZUyEMQ4dBz/
MGMttexx1SiDYKKQlkE=
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fgpwv2Gv/bZA/BQ8dxV6C0qsEHWt60NIacuLIivkM16KKN1kvdhzOepIkp3uv0yv8H1uAb3O6P6r
OOi6Eyy+5KXqCdj2Xs22rZRfcTZAgkDFkNhCT29YHTCjsRIlLXv90nKJbd5icDbxVVE3BiiXww+J
G7dLCmBkMSn1c0mY4vNLQvW3BPio3jnvd5f2db1oOIFmUVCca5jjB+VBmIL5nOZdgFtUV7X5ovYa
8UUxcWF3rMa5aXbNGbfOjjiITXWr2W0x6HN+AtxEh1R7m3n39uSuUtImoyWFt5TlqHENNmLMks1h
1xzJQkKU3QOJfM532o9wQWksTuiQgBx0BgHGUA==
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 36624)
`protect data_block
upLAU/NTr09rnsiJI7cKuGofYTvusH3PU54RE5/x1U+k9ieBnH+scrHOuyyvK74ezQkXZBYVGU/B
ZjjIQfTVZMir7QYDhX5jADZj7UatJDyJo48s8TC0b1j9n5dhCaD1wbpQQbU1IGekOcRYneC3E4sx
n9UsjuM9F9fSVgqBzUE8XHIKMGgO1oZk66/YOtqigBZm3fO+GT9gfv3XhxIUGXMqwlxMm+wj5Y/1
dFo3xXBxHa4hnikUyCdWYyowPWQIyyuH0hEXpfYzRCyuJTLut3g92fbkKAsTvMFqdWvrx+YglF5C
j7r4rfR562h/CNwnmIPmH6hYNURG8/nlUywRSnDwGX2J54MHbwAG5vG0EZNVT9Z9Nq0AQtA4wyVU
WopKgxYpN3yaA+31p81n7ay/+JQdlcWb8Mu3z6WGJZKW4foVwHaoQ5t1A0c8hIsZVL6j53r5gewN
0E0e1xLEXhVSN5EDfYFzmnfYVR/b6yl0FBoCvU6MXfyeZGdIZGhKZ9IUDvQZ3GYsVVX4cuRiqzkA
UuI1BN4OaE4QnZ0JmKYYf2zOjKx2dHTIuRjuyiyFNzPCNkyAhRvx7DwR9Cb+q7SMNUGiI4sPrTAF
DgDjXan/wiUu3MuJZWSlrJkAgBV8HVOLqjQV2Yyyf6KKJDuK0oV/bPklWR4TxVYBJFfEtfyftBr5
qcT1J7ePqMqdUpy/rZBwJ13MgFwLSWg4koZCvdRFL2hkomLbQS4RRvppPPNof0/UNQX4eR6KbV8K
HuzJNZKrDJKZOdBvg5RrY4Ih4jl9DO3VTFyL37H4ow6Ye5gEZDmSeNC+hNaTcrXLHwOrmUKX1kVt
udiL0XKGnTZYz/5M1zQHG0JCAwutyfaRtwjd7haAz4nsR2kXnNVKDhpQGHOk8XuvkYUishKJ55Fp
OYzGpwkHCUDFDK2yDOYa4Ds6ZNRJj3IozBVPuLYAKxYBXgcgWjeOx5jRdcw0L30ZeSPSIDp1/2Cq
Qfd19s8cUcK6/CxZQ9GD34lT17WLCPDy/HIvkioXgxgLlasuCUKRcW2s2ZpeePYDw615EGkWskPw
nw0J5o3HZevN4L9inWUaeEh2t83IQITdJPluhl9C9IUgxu1+6aVerQNze4GZcw4vdrsA2q11RJs6
RJWApGaNe0cCedRj4b/qS8XsnrdFS3z9DBQ3h5jnCldZQn/B4kROlGjNRwunEN9rZ/TtXnXl4617
PNB38K+mePxI0PLcYWb3FGVjnUXuiDT2KSthawRJWz1+VIkn5n4D/91r0R4cML16Ey42gl7wmOY7
N8SGOknkBtvMSuKEXGzQIkpkkGHirVT/czL5bMmiJe/GYtUB1tp/z8a3wXHVuGstFbZLriv7U5E1
hnavkrshgWmdDRZWkWC1tOdvDZvfzqsP/ME0aTEw0Wo3VDY3zP+qZfmNshMt9cp7R5+WIjWqk13y
5pEkyj+r866vl4IlAVoOteoDq4a3rr7+UQRfy38vTJmoKx5DG9sR+36jIqQbPv/36S1Kxw4ihk4v
IuVJgC/ZpmRUL9/Ta0wh4N81eRpCTwjJX2lu7xw6MaW30uRvAAMHV4OAO9GgWqV3Xi4u3kD3181B
qJzlemN7oOF0Un/X73jnI13L/K7rkC0lMJWsDCHEi6ubAR6nFM2hSjVElSswSdqKYn4rF3RhGAa4
xFS61HkXkEYoZ7cx9meN1qjF0sEv1xHJRusbMm5gTV+7uFFrUxpHWRKuPZTlmcUvpm7IUIoO1DDy
mVV/ECo+S2/qBtzA2yXbZqwdoxPuSl9A4llkaxngRhp0w8jKhSI28bRBwYWgTArs+GvRglZCGxcX
tPNWzhEfOyA6JiSJoZf2EcqzJMil11gdKy4pSVTmcsFV37PAotdkdYRaYZMTvaSZNO+bvcNFroT4
cQ0BH4E2I/yShukNvE1HAjqtB+/5WCd7+xeUfRmvfSg7qgKk3Be6FgAMLSAfLXnXMC74Y+gwj7HC
Vz6y0pahYOl8pY8k2+uNw4tYebUqcWmI7N6QuExUKootPdcriULh3bex9lntFcM9DmwLPTn/htOz
fUNFWVggsj6vHTvNUKhZnXd6fWOcPqK3ZMPwX8E27GOQjbUuZyt8hpPD2rdOsG9MC/ugrf4U/x9f
aIJxXL3VS+faUgETprnUEzPEMs2GUV4WFc2jvinOur48d8/Fo9/YyrZ7hWC0zprEU7ZcKk7ixR2K
gOWQqPRfQ8oKpQliPNRJNIpJHMIMif6+ZaKY58UXbqfihFd9b3ZxhbvG6Q6T3/K/4qkkCQlcCOgR
sYw47n9smx03ZAIeY1U2fqq7HSbrR6QJ4JyF1MraVEYehH396y2pEN7r9XU36d1ronRgjzJDau4E
6PpSqWLC2TIFTI7R09S4TAu32pdsT4pyZGsnx1OeBeJtlBT3Hi3IyNZaniyCF3dx4IYZaK3Kl8Fr
iwrEry5jsoC6hZ3SWFUEcHpR4xVbsww07Gn4W+FvXxPKEEoZaJdhT4+emRLX3V4WTfKDxm4fHdQb
lU5u2BDRpzgDGl7OiPcLDzg0C/QPlmCKYX9DH4UQcU4EQ33hnbvGABL1cp7+un/LzftWJd7fT9yB
Nqs1YQogxBdBubRIZwhs2ma2TWdTr2EXOVj9fcBvXFInRwV5USssbrcR/5lLQdokT/n/s1SAsiU/
0gG2WJgS8HHsnuPevkQlIYIUydaHr+IjkKERL0l0xY/HuTDppExzynOQNEm2gogoAizb4KrQDPoZ
08TTHZ4rHLwManwqBRgOhACpd0qZ9HRig8n8G6r9Rteqx9OZBYClDJiQ0bRPV3xOEo6frYY/9gTd
MkdX4Gy2Y4bYhuP0mAur/JFES8n/bLLIwnQp84KNXDRSrdvZefP2OGOfSDAzvQUp2EOw6/Ytb/tI
e18C/M4nv87dgKJ4luPLjID3MNAxr5vEpYeexDndS7KzU8/MGkeOhdgVO6NUMZsVIPc9LUtFDidj
mevZ0dqPp95rHR3xb5V8A+KzeUrneLmQbi1FwoKS8mhc1qbLs3Wu7dTlAp2ol28ASWqembZju+Q5
pTd4uTaikObexIRtTh51re5skXGPdCjgeAtf3oSTOBJPj1v/ejc2O+xGwM2DTVPmRCjZvtwceNxB
c2cCJJG28/4XelpC3FXC01kXP/TuP+Nh0CjTE9a3ro7SmHsTcL0rm9N3g2+fE1+HVFPh63HTsYiA
XtjvxJdBKrYdony7tJ1LBz6Rx4vF+Np8EK0fkLnxBtCNzVxcP/jNC+Ex/RW5bXN164Tm0qdvotSi
TK1zEGSCQDOLTkwfADvhI9CJZk24D3DHp1Nf23zAmfv1fBR1QLPA09I++GjjLxQu/iT+O0JQpljA
5tlkeP+KfZ2yRlodRdbb9RBL3fES19agdRdG0CxXPdR+CmPOk2QCXlP2M7PQ8/l1exxjyw8b756S
z0UY3ouGNI7H338mmYKehlyJs0yugwa/5G97hU+lR8NAvxbJRHXKXaLRUSx+beztgsVQY7CL/inO
M4erb+Dp6bgXFtpxudFTXSEgf5ePeaIMKU4QF8H1Szejub9yWvBiWCqkk2cZ7zSHnwrQbFCfox3F
0ILqljXc8dQLKTZ0rJdGjQdwcUpvpe5oP+RpWw22u6cMqs2V2v6lbReePOnAQLQuSGWTyARDkKgv
liBji4D0uAF93v/F6ZZDaehE6JwMd6dIaxm4emDRfOF8GLqiddtTCT/SimsQr+uLc2aHkt7biDHR
+NJP2NWXhHTH8Hpit8LultR/MB+9AuUhXngYGbNZf2go/dluL1IX9zRAJe/onXxRRKyNb6qjC6Sg
bqxCC+Yw3YpibLTWM4GGuiZ9DDd+G0yN6C/DiOko5RcPCnUmx1SaPqwqAuXYwvo3vepcO+6+YGWF
WsXyc/Bo3400YVHhtFAvpDGTv3Ffl7YBT89sjdfU2j9FWm4ni1nYok1Iil/TYROnOoez8rHA/XKN
pRg4rx4ANrWYhO/TUBpX2tEtjCa/lxbJIp3V1EnVBxHxfkGPkDjEXiG1d/c1Jjsxy4P3IYiMlVt5
1cI6UNCSatgO4gXTmN60AsS+obknP4KbjM36/k3a9jYttSkN3LEGEbcf4T91AyzKRLXrP7J7e70u
QXwh7NB8m3ld4IauYRzng6LHsADBKbbooIJm633ydd6Z6YIQbnkey9FBrIMKpuTaldpljSo2Mx8x
PNcxsKr82zdQKMaUDC1wqw7biop2WQVq92Ie+WqW7XjaI29ChACirZdKR45dDIv73csIMlLzC/iI
qlqxG2KxmhqJi6Tvj5nZY0Cbfdch8KHDdsmuwpcwGntgHTq3+zezYbTQbThccCIMED3btAnh10vy
qwKoo80+fTpY6TDWAuB20IzEUTmvT99Skh/5oBhUkQfp5n1hqqfv9fR/yqoHskQwem+3R2e7RoP9
TWxxhYfDR8tLkcXn1lAIjgK8awYae/C2PCp+bvna0ShukOwJ2zw4mcuMNMU9BRpXjbzz/QZmkwfu
j1dcoQ6IAJDPO+F21V7RNtgDQ2MUZUCWwpc8cpwpxcIiSpga15Xb7ii8Xw+h3438/MgwBytgtd+J
ydKeljxrPR3OiIVGCCxDdT5wtp2uHZzsHk/ug4/WxnAcflz+fyD6THFoR0xWv1PZ2CYhIhrJaEYr
/V0X5LycdBzS2J8PxEhy9aO9I9oHgrsD8Mr+H/DxbTpKqjyf9lTMHljyN/bHr1SmU1G6yAZOEOwK
OSAPrUvAcQK4kV5AEKM91YXlIcTczsHfADuAWIYpzB6His+1KRAervwxElnB4RKlRkRMDqr+G5dt
2MOu6mVbEx2Yg6anJBZ4vWFoyOFLetJQH1d2u7x8srTnSNOS9/xZl16i+TLCW2wx2uHkSo6WnuUn
XN66EdH1V9+Q0vIWXhVjaF8OWTB4CaufS/ACnYMXpM2owJ+ncy2H6fj3LgFgxuoceD76cNIrFVYF
MEwZkLU85GWl4lolzk9LuQ3RmKzbYtQ0/Q/4UPezV0UmIeCVQLIhqjRztcdTUkZq6q1ob4NfKIkk
4aYsmUn125zEUYOkBeVzsIKCBuasSFbuzSeDJsjnqILsky2NZ8//Ay+VoQ2oVJ+FuAWcezqoiDeA
c6E23Ooed6Ywg7AXkL7ayCj8BidXw0s+FW0CeYi5pOxLRfI1T9RQxarHGzLomwsfP7LL+G4ouIza
tACOqWQhBIde1o34Q1BHTXmXLDMZWEo1bxn9dEfj/LNo8dWmCOSurrxrdNRbMFO891BnlP0lEnbj
Ojtr/oQkmGXGve8QtWNuRtM0NqwwK/dnLEpqt+xaEgv57QTzIjX3ccaBIVJ0phKjYRTGScxFKvv5
j57mN4pAuxmOXhYxOGFEDQnsixe+3A7c8JZZxGhrELqRwQsoJxgsnkjhTghhCx308Vo8KnqQHSvK
55ie7zLAwQiwuzTs5Og4OboukpeVlzQRDiHi489op7Ai6IxDujig3sqW2i5MvQC8XHrLRtTXCPo0
4+8CsXQh23MjqrWvNJLzID0wnnNDtmeYafaQYWrClcwaGOM3M/A+wHOKOFgBgs+2CK9+ChBrjyKs
KlraI4eCLnW2/F254/LNWrpGykrHw16f9hqJVd+FoCYMfv5JGvjjbCym1oNtDg7cXpsnFGEpN8Gi
iqEurnqaYhMtWXENsNNgI5IEbp5ccoEqpDYstBLV1PFZHiiQ2pSy0RceDeVzGlh99nvUFY4r9VER
KPzKhetofIVYt5VlPrfjLydYQrCwQMpBETvkSTmKpGx2GkDO0IMeCAEiKNOKvc72HSJUodfjfGA+
24O0eAgORexEQpuM9pWMMXyR4Pe0UrW1oh2IeL40qvz8crYKzxg+FknFA5LPS4lemrxs6/iiJ8zJ
YMWwJBVj38al3KKiG31GZaHRp4WliQWxXAwLjpUiQ95HegpOEday2WmLxA6RUEUrMRDIGzgOfpao
YnQ1h3ibpONQz5CFuQ1zHuqkTKKQ36QzmXLPoXt2WcjD/XQ8Xp4eWGq4rQ0CMF47ptY5eAWeqdeH
JFAXsTvVXyHfqufuZQ81j61FG2Bt/ATCNDwZ0LwwPmB2/Nnh82l2JsuN+Oq43mN0wofaWu//IENK
2S2EBcv9p/y1sAKKE2jvaQYO/+uIDmKiiyGHwdVaUOBy+ok1Pfz6i3bZY1rYLB5g78hwN5insCXQ
pryK/KvjRRjh572gmpgx1GUe8NcN1p8tJgBv3srkfpuyJnKam9Jgv+ZLLKh2M7y87boKNBlU66av
eBDq6XbCD2YUjy+2Y6z3SojLGqFHnumJ6SUuxuN5b9cTkj29pekPcea0bgAM/meq5shNZEFyUJIE
rtCBNIlaSc7bjIYgCxWUqsaoG9HuUwlEvOHoACmXv2yJJqWbbgUhOIWv/Ui7ayYGy5CM1ysTMRA9
1SSTBXiQTydpBYEahNS5npucjfOOg8QCp31z165N6f9w7Y3IPFLeBCB491IQj9K7JA3HHVN4B3E4
AJUIZDgGWVj5g1o1VmRsbu5tVP23o+nWzuzTFehG8PP2XYUIJaas3Nl2IK02G6TtEBIhnqLVd32z
+o92KADFnLEQ4jG+JYLlyTEq/cNq71euIkCjfIzcAudAtWJZ9KaNMzOU6n1SudZVTSLsBhXrUlFr
GfZjl1MBrZPYE5i+DLRBMGKZwgBdrhsURePWbpRpYFa09+1X9QQ3yz48unht/bFGgAtLYLrf34sN
f9pdTU0bKgIwLkXVvGDt5bUlLWj5Ky1u0/SoVt3zzrm5DAWqxDoHElf+pGPNZiFofUn+xivFb/ay
NOfsi3Iq6ztdNxg9Ps2PELk9ffa51Ant0oY5h7lNdFHJwlaTGGb2MFA7dU51Sn2Uo50F1M0fbe3i
aWuiSanHcgUHVaCClqBlw9wtNbYJ19j8/XikVGc2Lp96JCXSjsFL6W7/rgNQrzg3Kp7r7bRv6BD2
e+U+MmAWBXLuhKmasfPNNN6sCrhg7O94odKNmF4JZMzqg2q4rbKFBtOXZNAaa60KxkRGkNSXeLTG
LsodZGWJefeVsKxwT5rMPFPyJFMJ4Wb2si+sZoo27h5hpEK3/EMV9zsH5dR1iSRbxtNszzJ6QVdc
ddr8/XRo1xFZ/kC/+iT1PnFHmCPrAlQupmD37N+7GRVmnfHeO4oFHoG/9HgnY38dHoS03DTdldCA
CW+re+epo9666zTycSA6njhHO1mDBN9Fit70rBKasl44GyZOc4pY0PJmTDBBoiUfAknxYQDg86X6
YFs+4pLqL4eBmmdSHFJYNN/yiRCF8vPZYM8oLcjqvBRC+N+T0oBvDm2xVvD7Ht+BrXyhYN3nYL3J
BdyTWYDRUdR4t9jEkD3TY/fYrPKOs5eZtw7L+4MCiAX30yLqj279AScyNLbQ3OBC+/h5NWejAXIb
1/UyVkAPlDaBbp5dcCyz9YeScH/6f/3qZx1M9GxbMym+U3fchNZjbgfVQTDjdtrXDBKSKe67GA3H
g3Kk3mZdTdA9DNzNuFLEEGNoMPMl4ZjEuwXYspShgSTEMv56gUhXvgdGhkNX4S/wytx5A76lXFdJ
Y3bGIJpycksKRGK1q6BWtvRJSt+yXwslbQHEJkdNdqoxrostv2n+6J4tIeYdK1vi401Fo6iyOf89
aTB7iq6Lw4hun+Rg6ADdGkdMXvAerQB3p6y5GQPgG4qF8Ou5qvV1jco+PAqYvJVV0U8MAcHmqtao
mOLs8T94slS4AEd7LkDBYJpANhYFXwXXwHsG7vJWhGByc2W2h5z3Vf+ddr+ZuJVl3qnlMjJLNk06
J71xdR0cgoL8vg5vIRjpUE2bS4cFYUe6qlWprLwhgXr/J3TpoJ50NC+ufEpm9fNqmeBu4/kd2php
PK1aIp4OeNz2s8/VBkjjc2SCmnvkCTHI6xjJJWeS6xPhlMQ9UhNbO+SDrdqj3WBtIKMgssMFbX1r
/cYFsDZcG9cJVorbFEJdR7Ky03u6C9emT4ycoMJ5+qD7An6XIncRI0S6IrOPp17zmqF6WH95/EtR
ibJJMtAU8pNh7xPJWEP91pOnQEvTXI1GdbDWNdv+x9b4CfQMUVAcv4K9h/n2kJE9a0G6ZZZ5NeB2
5femg/sFWwNoHVRFeIjocbfF6+JzkEYAcADiDHUuo8UoivjI7/c9pXp4KzJo/Yr3AMVxbP9YnyoM
sLBuxQYsZ5IWGlva81BIACguHWn0AY5ign4CVubXEpDUUvA6AmxXVXzmKgfOpxvggKnH5PMnu6JJ
klNZWmwgtudpeRtutpMza1goxkDNc6+BTT3JVTIzZ6Lv50ohN/uutJyh/342vTuutb6VCoM9RSpN
z2HqzURZCc3TWfJz3U+Kgljlkw+ZOLjiNMfkWhz6QxIpnQOB466HW/X5w9vjvn6pXi1ksQEBSdAZ
h1hAS5yOS+0k7RSHQd0oGW5MGrzReCj/SSp81RezMz6IaqjnYiDhzx6t2kWcgjR1ed12DeOvzfLz
DPb8oBGbZJooiShHwUU06bs44TgRt3Iep8vYHNS8Y6zQFdRcrRu3dIvuLmuiPNk0ScMefT3l5mtA
iwMbJtoOO8q0HPj9nxu1Wkc8SEXaYA3xD7UOsMZC8pGjEnZyWiGv3vvjhh6Eoyop/pGDIE8/BfNS
ZlB2Jfkg0jQs6Q0UkXIGSmu0zasvmLPZyD/iy+ZIkXi201gu2ZPt1HRDIv2asnxTtkSWZK88Jeat
PSPbFU3ZkqOE/timVAEJD89exx4LbnfRs8M1WZAxkHYCcgXGblmEwwjcYPIDGL9jn2kWodbPA2AW
mUmmkCnA2rSQITfvRWsnJ2AkKZaMJO9wuQKZK0YF1ho7kID14BM7NTjq5gwrwv6SU0sCa8glNHbR
QIWw7jKXK1d9G8d1n009ofjFYbx46627x2w+a7e6evSBSyh0U22Wx1OVIx6NVVAxORZWkxAMSdrH
T52H0GvzRA9WxTf9tHbBcQ55LwFUlNu8kX2lFOehptzFnm0AszaWNgOE97i7Bp2QJcYRL9D+uxKr
vCp3h6/37ZL2RohNYcAjofyu7U2xa3nUNe9AjYFKuSe9g9qtOpBZ1TSkvQZryNzW3fYVm0qtLbm0
h4nit23oyB54L8MT0R7/hP8fJwJq4C5H2E62WikpP2OjLO4DG/6x3tHHcS/q+5rZyuqI/5Ox4LSp
2CrUw6wzwli52+iwvQBh9QvT4H4IVHuCGd72EoravN0iCWv5ghViek93qwu+19PcNXs6zhCkl56b
RAGo2Pgh7wear5l/Der7K5qYloyMKuXYpFg8BrgE+kGkin4HdjtKCZbC1EfAFccxEN1GaqhfYoZG
jvtcB8k5QWybNUaW/7DKUzFY8iP8C17PO89GGGhbjui5qMg+LQF9DhrxF0LvA9uQtBgCU8sxQhP6
ujR4QPnDVvwfXtvnkVN6V+WsCkvoUxf4pFTjqnR+2YQ3bTmeqjfib9Ux9hJIkZGMnt5GYpCQiUF2
aVt+U1Op+YMD3FsDzfpgMs+s/tPBUponC8qmC/wRDDJRlWXCl/Ug1mnV/v9IjvfBuiZlNHVsp6cv
Jn+IXF2FMt13hYZLfZRDESkLnG73XWgaASS7VpqSFf/CXbIyxWD4gw5pwRlBNj+H/ed9JpLuWDeZ
dyQGjudWs/X2/TPzd0xX1ofq5KczwyNCXzVSyEBuz1mZp7UG+DfKze8OFap6tWEy9L0GG1zSZftU
z+BXmjDY6oq/T05mc2vchwJbpAJvkKaGH2ftVqDzm2oo/Ry90ONlk/noaMP8kf/EwwrgZgf9h39o
PYP0i+3GqERjBd2SRuAKFwgPTXEyeOLaPFzzwXAKHUZ+iyHl94FgYvMHOPL+tCDyufO/MyKamBej
3H5rKQQTi80SRg4Yj+LC4PczOc7IsK5AN60Ff/7QkQkQUmwDAoRaEzeuHB9TWbFD2Alu80PkWw+j
sz8nwPzhzb7EarFVOr00wxp4Kty6LiZCym2a+yqa0KmTynRKH9DpQIvoadvVwSsf+5Qd78MBl4zv
jhjEl8im+WxUNsLKK6r2ZYaq596eirJUO0V+5g7GcvQXcXY3mYLBmLKhJrn2aVw0YUlHRd+PNLHf
SAkZOdXfAGIcNVNh9CP/s8UDU7kjKXQMOYOxqcIZMKIxM6iF1rsFX+hxRjlbZ6CV068diXv2NJ/E
0/quZLoTb/jGj+7YTVDVusLkUuNcMxZn2cKaRtrEwQ4gc+C6QgJiMDacOy6CIfim3wEvoN/JV/jK
EC76uFUGpagUBxRZlsCFvbw4yeJhmaQGXY5dC1E5rRCz+zUQ6+k57Kp7cqT5TPhZx04Cw/FaMo7C
5Q8O2H9neLbxrbZwIk/jnEeJSoWPs82gJmQrhyNheERK0OHo9UMh0HM385082Xg9arWaLbOuMO3R
k2EoeGSYfhCWwZ8/T/EK9dGVdnweUlOL2twgvslneQLvEuNzB5FF5Zi+pbESwwwlXtc1hb+RyCuS
rjTjHVKvM9PIrO2jmUgMODXolgI61VUF+R8dgU1EJz9QkF6+3GDlqzsZ45ymD/9k/Sx4yltw8hiI
FkAbugo6Y4S1a/DR6TNjH80B/V9Fcob9cp2qJhwHdCoq92P1Lw+abTBPJHQfbhfjPUs5LowHVYVx
2fYmqURGmHytQkq3edfnwxzhLxaEjP9dR2W4i6/HnVtqABxUtptUQB/z72kDmCxa5QpBMY/sXmEX
nRdY1bMZjY5wQw+r5fYosYnAg6zVhFgDVPzsksFaFkHWVINl/BmODcduysw0Q+/mMyxrJweNh6C1
j9Dk/kPIFX8eYQrFR8GxB/wLUsloz3BkXl5WszJUDmM6WHl6ZjA0ecXlJI5lidzy5tqx+YNKo8os
wKfc0MVpciSlP48OgjpmkwfVCN7JxFU/QRR8S3oqYzm5rUizl/SY0sArNN6O9QDY7y+C11habE2U
rYY1af67PEAEyYhoT4IQiA211XUN1A6KqIzP9K2M/0aoWWDH7BRUlOdcS5LgOyKTOkMHiCLtvaBe
ylViTCd3EJARhF70gdDcNZALKY6vizsI32/Mhr1L6N8s17n4KLSiTpgR9wkWMiBrLBXUu6za5mMF
pU1ip4j/IEeqCk3InHLWv3U2CT/bx7FBomU8kMCoh1tKMpuWV+H88VfRxbHX0JIaIODuMdTtqD+o
NX+ehrN0gzxxrvBBGZu2s7e9rbsOIWGdgH7ZXwULG5P42OIV0beVjSY5mGq3BA1iPTyFBh3xE2r4
bmxQoEGgSpp+W6elwpH0wQMvZ6k8uOSBq0ReWIzmq80XwNdFgJoS7PscnFgTG2PMm2cZvzFVJpcz
TMkQl4mZa6bzoyKljJWFbNJ8n1i/bjxmRPFOAFPY+e2q47z2A8VFtR3XQlSSB46CpYo7ja+JO7v1
EWqu1sqZKlLYwty3ewwt8rg03mnO6uWzWLlCIO8b0jJLncCwMwUrned5iz36nzEd3gtkzfO7jUcY
oQAFeLi1dqpn+MJSX78mEylgtYw7/R8wa62A3kZhaP4TytSVDzY7PVEXzFiPt0cYJTBWE8L2wikb
d1lOOghS0Xe4fvwW68AeEliAI2FCYRh4YUKBsrNDxVeAg3rkov4VebUR/tlp9QbqOSOHTbqhAr9b
suVDDyBKD+XBglRHAPN/RVEITqeY1MglqfgAWPQI2NJfJHYMQbh4eg9uO0NWSNZem3ZxqXOHKvzP
y88c0bC2jfMNA4qxqkkhZ/jenvm+MkNzYpcrSU24+S7RW410U9YfA0z4G/lplC6/66ZdkeEQ/7HN
G9W+PKt9F6uGEGdm/e7RbUBzMK+0vrVZcp3cnJzITrURZRNqRWonhgsaBlDcwf9sOMUbdSS91aTe
LKpxkjX0FPEzsGioVaYcX9+D03lc0/UBKCwwrajjbPKqv/qnlOixQh963ClbXHKyCNkWOgdA0KcJ
eSvehVInAhodSLEaKVVEPnbPaWnVrDaEuj9vX7w/g9SPT+STIX8snSMxjnkstd1Kv6Y4rb9q8lgj
qe+LTgGgwabpzwF+AGz7STN+pIdvpYPqTSyuusbEfIfrPjttadAxSh8KmfRREhb1wummhthGUz/8
+VXQk1emK7mcXD7SI4GsE1k+p3H9eGMQ95guryfG23NQshn1dzNppPcoLQxMjfdXi5xGZWadsU6a
oUGLWEKe7zbZAkT3R67ki5XiYbgGUj5rRMxOb/3iploilREQpRTnkWmzHce0deFNVXdV48s76oiA
1wAMbD+O2SmOCtYv7CbS/z/58rKpcfZC/b5ynSwbldj6t/x+uwViVqAVJghrTfsH1NIRPvUJ2RV5
qYO6KWPTRAReAQvGZLuk7iR/nD0YLrGLq1i/FuiDEQGqyRLgbzWFQqfDr7sOWz1C4A11x6Q6++7y
mEYg6VMMcnGBjE5+A+0k0TqPaU45GWIFF5unCUnPSQsdD3gCX/iT3vZ6lBDLA9lFOwLl6TVFgpOU
dXJWZl8FbvmLV6yn235HDeIbf1stugsct2/CSWG3NulbmuzMf24WCGfFUREETesNwMPbJR6Dc6kt
qvRacgYvlHFmted89/viLuLvJ2RQtKkwLSuDsL2fEr4GNiIXVCOi5TWJiC+RZ4tv5WisyXMczq7H
kx8cqRs83KrD4YBJ+sBmyXC/mDQaRsKZybcf46hl5+gE31l5CzqkNTEDLpx61BVAVPm/e04eCFab
aO3Gnw9kVWDc0xpsPpOL934wG3kfrwzOcb3Bh+4wo/T9Et76ewdhYZVPhR4qIKP5SYuPHZ13IE7u
OEySN/UVQTWJ2k6xkc7knZRj4vTh71p41L7sxjVHaWAX9yGuqv4BK4L/PqtEuSLtCpdhF6dG8ML/
sNlxmDDIFDUuu1cJg0a/hb4mIYI6HCZhi5msfbffyX9NGIjkZpYvLr0C/R3tHIcweBeMAsLBZ3lp
54FHdz802gqeBdB7u1xaPt/lXrNd80bOTLbWyV82Z8RYDpBX3L4MR1A9BLzWCRqk/Ad6Jmn3KGT4
9m4Pb4HQEEp5Bwj/+kDfyAoWdgDoTEHLYlAFnSIoi7f0mFk2ojEyVTu7Pkdp+C6yg2J7VE8r7+VR
la9WkQ0Hk/RpoG7p6NGU1uC/lJ5PsgJOMjrP2xIVE5HCYN1Fj+hKY+NjY7t6VPwwf68qqWjd84zQ
CakIWrTTVroINmK4XjL8uSihWFL9vBVRkgNfHuEIFnRUUASHjSGLd+cd8LH/xeAqWMG+6klB3NOV
oTqCZVx6bqse9xCOK0lKVWDYIaL9ry2/c5jUdnz7+gszsHIxtJ94zEOV+G3uHqVHp9FLOTlED1fD
7O4yCMvOwQF51PFP+AOeZlssHRCsnxihAf4VgFaiz5+AERhkISdsaS4Mo62q3Jq2O9DCtMKYv81O
AHWM4Q/dQUjUIc3eSWGYW3dTmyqYPJIpbZmbBd73LWmOsaRVc36Fxr/9ydiEuvuyXDy/1WpRpkI2
7Vln4b58PlN3lp0rTt0Bu7xFjfs1/Z+hApiOxiG8mCzABjMk1f7CPKAB4tP3YOuoyXIBWx9kbwC4
Aa9A9qVv0T2D49q/Nr+VthlAMF2ex9Nd8h/COot1ORCVStR5vByt3+MAABOFxUYCyB3ujV+AJID3
ccmOMEtDM2vhR7nCjt5nu6wURFEA6mxrDAmC14UpLmzlmpJA/4JOJhQEca363HlU0E//pQEzXmTm
ryqHkfpuYRU+ujgG79OwNnTP9IdCMIOFpA694ILbMT7P0VAEgmQyFFed0arUD5Ox2n9ZVgvGMkiI
ujqqea7RpPeJQ3ed3/8klhKq+3sZcTUviI65y2DCnvQB7fcP+/dhCvMHitG56baJ9f08nYXXCnZv
0eLrwta9Ia0zd1xBbN9LkzDs85AjX+bhOLco1v1BxbDScgSPI9+enXnQZJJYsq75heEEhUYktsza
rpcemrBKotCOD0ChdKh5gTbTJOzHNK8PEFik5PDRsFXooe0IIHXc8mPNsrTiMKRZFV0aNMBMrp3S
FBP2ItcQ9Ij4fO2ZfJUu5D6AxPktunOow3IMT3GpOUSmLEvKJ71aFiSmJWm8CZy64dIINtCPu23W
BGQnoz4r643iYxuLJka6LCIwSWqlzFRcg7eISAUnCDw0eVKmobtCMCsKYYfwSd6466Hl5XF5hFgy
gs5tvvviGL5/mTsPw4BXYvJh6M/bogj8asAMbmFYyNzpGjvHMBVWZF2RBhVzujZb6qGUf9Qz8XGU
oLw+efIvZ087UyrDHoCVr6zx3wlr1W0UvrYZN6U3BGXFywM1Xgl7K6vKFiR1hL8wNsGUhSxR+vtg
4+ckHFn2wh4BstTlUTJj55tlXUz80ZOy2MCUPFXiFQ3Q7LtwIdmY87jn1l1jwCaqf9Sjzdu0QRZ+
AT7MdQTr2WUJ/AdNLk5SKtaOKcBtilAZw/fgph0RmQmb8vqIclwRaTxbZt9BtbjEpECIEEXQ3u1x
hFrkAcAfw1P97rhtzMdZQFg25yGH2hBE+ZvW9y7JR95vA5V3JqueVRWDFIjdd0sUuaODqCehFhWO
Drq8hZcpIZImCfbIJmLPOSXwY/gjFHpKeC+44DOw1uGcPayb4QuCEQ3NuoZVwCELxTIlWDA72ICt
0dPLJW1zbGG3DwNO0sdoV+jXZa/58aufwGJZUMDaV6D598GPmgK9qIKgaKwFKKi/0+/sGhBTUgcj
YQ/+XcyqhugS1Y696Hi/bS47MSq5AFDibGXT3QHUpbB0AJxNwsNudCg7I3PTlMwKHv0LTb7E03V3
MO+wk4deHyX1qVe1X70N6z38kShCnSE8U/gLKF/0donaynCvLtEeFCzNXDrnqqI7ly+savxOBtWG
PPA+19Abnq9ME+4CFVNvsNTVPOXq4yfuks0IWUifpVYk/S7WuoJVNU7+UsMXntwauyS5ZvGxwOnF
SW3QCbLacn8dqNaRoS+31sT6iFtNqEyXORRxoL+km6SUDm/md6cySqrUi6vYItqcZ4g7llZ5HWQN
TX4zc6gcm7oqg+uvumukC0XUNbhEXgFZ78AH7ODSaDEzFSXxKzy8Gdvrt42X8DQB13b8+GMUi5pR
Z70qPRo+8UM+51/k7G+7WYFhY/X5UOlOcXRTF2JV+6krTRL8Idwo/7bk6kUTzKxyywJu9Zeu+IdD
DVXPEYXUBXJCaeNl87NCj1eeHQ+XhA3OZanvhJf6a8xuS9BGwiGFwE3Ov52AKPHe968RCwUDYWBH
Z0JAYTk6uNyzy3DQbFnsK8iwEAHrPV2OPXmunRzTg4CiIfvC86wAGZWK+crZX50glywekrUHIWRk
hOFvqJsEbyOtNAjtNOv3g62AKtoCnmXrBafqNkikEVKxgY7r3N6HYnsgxzXnkslERg5+l+NDE/qc
sDBe90ViMqeQCHQ9w4mY7tnzFSyE8NjUdJ6NDob1gA8PKk5KodgG/5+NNaO/9Ft3rwI5VOGL2okx
e3jmOXVYRDPLB0i954Y7z+Lk15BaZLyURWLQ5YcoSBCV+FobDUdeFlLTm/mct1uegx1ohKjgml0i
xxI9yl1yYqHWk2PPH27mWUdWwQfEh55wtblu7B253YIlzDC+/6XBWLuNSLpFMr8nn0K33Cfi9eGT
NAf604LA63kLPQMfsXaUrbBgUU299Y6hEgcHJ6vSOBvdzXpsHgn/sphkaR9mVG4jAr5T3iMFirjB
9B85DzlPzBdM7wMOcqPQT7671om7VMrN5G3GPtHaRRYuPcB+QdhQ7IdAElGmu3RKKEBLd1vYlWQF
RoHOoVsBs7zgKflOQdHJ4qorMJeZ8labOQaLI74LIYFJQ8yQRxdes5fgUdraWx2bqq1KpJBvsBCP
h+5jMGRGredzjMzhBKtnd34cE84a7usCN5E/SKLAN0OmBVl/klX/jj7FKVxUtUAP48mts96A5HEG
4FeStYo41i7Np7tOPJ3ZRwle8ATRNPhLjWNK3Mcp1GIqga+RY1DPvL4ZaltonfC1kwDhK/SxMf1a
dfdo5wCd1ZlYGs3Jxn64z2NzvkB3rlMNZ8/zJoqgNb3jeAWcoi/tIUXneFy3iNN671eDlvSIJt1t
nP2UgEWLEK2RuFwD/3+3sVxA9sxAEcFzuRdThIVxeM72qmSKLXIOMGXgXKpATDKf3oKxi1vBSLpB
axpDsJeLZ9I0IJohXKX9MVE39xWTr/EmVoMwxo0uLoQgJbQLP7BZvrHIIMPH2cEaw5n80za+O260
WR+u/IHl8FAlqmwBi6c1odAQKPxFwbDPtHIu5hEBWmPdMKW7fAbQHc3e/9ENZ1Yx3skOn0FqHLTQ
sC4Qt56mdPA3MyoE/TU0Y/6rHZUaF1eXnQSk2PmvqzzO23JaZfDCE3kEuv42yd2bBsJ9nckP4wSc
dyR36TPLXnQKTfPlwjbeEctF5u5HM81qOVrI4KJ4kvCxvAdxHs+gCbvbThVWyjK+OaxuJa7cUlpn
1kO+AllMOBm6CZn2ksOApFe0QZjMSruwB3hfF5ZLmS/bgPz5+Z8mnrSgkw3F02uKM5oR7QEwl8/P
Ul/Jz1SGyQeLAsjL40nHUQhjsCCrGW4US/P310ocyVTOwLHkh+HBOgnriiZgJAPjOc6UQzfR8G0/
KNfYa/e5Bf+6KGNA7/pSh6u6qJAOsUdTacM75M4lI9LGeAnu6CaPDg2fDtTQ4nw24Pn+lItkSX0M
EjCtyl6KUBUdtwBnA/GRrzkPMEsjxMFBJtIjQBXF1Et++ktyV3B4blRKogHlZGo9tJX9iuW9yZjo
2cFKQbt/mtuPbljpGaDHLRwTrAY6fuR7QWSG5a71HHaAjP04ZLxnRsPA1ckHbkV0Vlwb2cuNbAId
MLUT2BPaZ5wJQC0ZyeKi3wgKOzlxL5zn7ml3x3JWI6z/6JpB9dpEaLjNZ6rFPxu7ydJ0gw+1zwMx
iEpprDOa9++ajotCTBx00YAEL7iknNBdChnVcOuRHEP+faUsfODXvxpwsHdUUf6Z21dLA7ANQyVL
cGDeyvnW3TK8C0oJsawpxtAMXVEUOh8hveDrqv0/x7+cPtk5pMaivpGTp36vgDYM51PyXgcTt1R/
UIIU6I2Ov8nRx2pA3PF021t9vGRxllSEMcsDU8Ptnq14kFU0P9cwH9/ruVUfROZmvxhpVQOvE3Th
yfXm+UpmcpXnk7sUBreEei0NXF2whMrpfs7SxGyW7FtggxsVt60KsHft7pozJ2798S0vTVmdr5/9
cXokZpbxYrc/xthSbO7bnDXbBWpHdc9jObDrvG4s5Ac8Kbra0kuUQE6oEESQ9Gpsr2v75wIf7L1Q
NK+bsmbcRhf3q54Fr0YTcTCLTbFJm+1mkogzHCAga+rvBAqDgEj7BD0yTz2OxE5QULWceW7+YCEf
Zgg4OsDJEhcWUFIiNwdeLFiSxJsSVocG8ds8kBr/QSpVEzGlaU+39TujGNmLK29Da80aDZFohbEW
pvML3IjcLixu01iMTiwawo37gcijQAX9UYna7ploIE8z1A8fHg5ECcuOiUbIPVFPf2G7Y7BwmH+w
taLd0T92RnVS5YGCTTPmNUtKNj4eSRI/GGlFsh1XOM6iDO+xveog06WfCvJFLh4jIeqmg9roN1oX
+AizlOOlzs7Xi07Q7YS8/zONZVqSWV9raIkkHIri2yP0eWzGWrRmjJ7XcAW7Q+qRF/JMwLBAhCEU
Uptp+7ZfWA9t8cjsoVYJaYnr1Cuvxj345kWeYmkYrcqKUsdMVz2Kd4hxdO4+BBuf6JaU8NxeuH/7
2HpmNjEzCJBPZxsRJRgIt3NEBxzbebisqGmBV8iJRIs04fHMfJPZDfWGM/mY608trQMJyCg4GFX4
/Tw3MNL0M0k2XRJ7qV+dADgiWJ7ONegHDxjHOraAbzO6zovlDh3/mk1Igjw2KZRJTgZcQR2dFIoZ
A5QszU/5FdF2nNM/XROi+ulqxqYq2gNgdHBvrblWQPWESXevOpHOSWuWGtrromnckdoUXOne+VOc
GYhujFQEYaXjnoJFnhezB0iaGq+9Oh4V3mQJFa5JDc3qTHbKsBrI38OAGZuGz6rqKGfMI5Qe/vPh
jVzN3d64SiBD1TUUoOo8JtdICZraqUyhniFg2D1i21i0PCcEmHVdoNDKioxbD4/oEahL4cKsPGkj
sFG8ckLbP+Q9xZ1RzT/KaMqnZsyzvBXj2qhAM9G1GpdUzJLpIoHDom1OQru3zRuNKZP+msBBVks+
dcza0oF/iyGjjZS5Yp+kx0lvHX/SVsElfFIK64FDmnd+RtNTWLaAZ/n18x8NCFRCWO1gbtPWZ6Il
32stsysPTC1sZejsDcaU+v1IxOI8wmXxqH2GjjFT5e3jmHbAGt/lKOg1JXRP/LtbRGdkwozzbZB1
FGvRAdnYV/tqegZBBNNAMIFrW+5VZVxDu+6cP3G7TOqUBgtjssokjSq93ikQFRnhIaRB6v4apKqO
zbCPN2r6xWEbG+6/b9hF1cEU0nuCG5A/2Bd8tpj5zEfoIimF5bn+FuMOe35+V00KVIuIfJ9hM/XQ
qLoaliv9+JMuiDh5ejTHC4M991rOiBjq3Cpal/Msm49PrSqwgjUbcduZGjJpXtmy2z9I0Jzh/4pL
eR9Mj/jsYDxumLP7DWTrTdjKhGESzJGVLlRVrGFdp/eWFHrLoB8nbvuIKF2zvukj0tfsVPog9LuO
ipTnIudkFqrftZyWrKfyvHKwbQJvVCASPBq/a26OZVYjhZ3+cMzg7/tFTgeOO/+l/MN1oJMmTZNG
ZvjD/2T5Qr7MFKsWNckxZZLrHL9Qjg8DqUPi1sprLIz1B+Z1DoZVF0mWp/p+7hH1+st3rxZ7ghr/
t4/b01VT5B6XDUQpTFyGPbMDEy3mzAIr7IWj6EMHEIj1NCeqSkmmJNaQ6NnIZa104iIs/NuKV5DR
YkzbxwWQTKR/0/JS2GqRXz2thmyq+qRl/6jk6MtdRStUBk9Pl0CUtk79Pbm7Jvh1H8YDHl+ks1es
0TvhzSeBYfxzCwLdUYRP1Dx2UDqZK+q5wIEXbwNuSD2ZczeA2pF/Eb9RfS90y9+sOBMzym7eui4h
OrxgKPGjReSeqpzStAV2QFXgf0pb+Akkc/CpuKzynphAHpbekj7mwrpGqbz5VzxINgurj/UC7uxD
Xa5iIv4JXPpb0I3cvA9DjkWUIWGvqRrkR7ElvbXb4u1LE90+IKKoBju6takr+b0cztlSg6yBE+bj
dvAVnKIGK6gaVMV6QJb2B/FGf5LhOTixmGNnHe5uOhFH3vVGxgwDKm/5EpLhlBsv4JatrDTx0FzZ
yQ+YGLL9qeap2S4ZmBYjWfE2kTYKw9MNArwtLdUCmLOsPzzKM5HY2hjfOWWwTs02gEvaWfDvNihY
5pMAE8QFEY9BsFL+NLPrZpJzlIF21LAKjOK00FTDai6mRqW446OYN4VVDry+Ps9Flh7qKQNTuyRJ
i2OuPHI3cLBN28/W+abLkt4lBgO6p+sbIfVAqW4vJQ1C94Qvww3rUWakwrilb4m8uC3WMu9jc6Aj
zgbcUIt2sIh9E3rVSIiISAH8rTEoJ3PxoOiF2wJ2votrBtNafY7w0kXj2G7u1a2WHFJI71qBRDOK
wFfSETx9LnCzRSw6ZG1Ty1XqiE8nZ0L7xvP8K8p6G/RKpLmpA8K5TwJLqVo0arpVL3Pt4DqjneNs
xO1pISxKzITPCoWkj6lvsiNU/Z5n61aiOhwe1xYDsYg+SWJtIhZKi9nFr7lN2z1l1RPuZhcpLtEB
FaQgTmmjaqVDKpX05fshwpit55Mf8pU4PPS/jQk3lBjkQ9INnkyUgYvD6Ifqd85DkEW45rrrghX4
whd0IYM98syc35fpc9vtTaGhAO0YJ1tgMLrqRkH+BJfjdziiarNhV1DHO+00WiIAjvxr6fYRDVks
OOpTG/QSP6/mMF52rr+t8kiZEilPZZdP13Sgx3Mh9NAk8Im1/XbucqR3ez1l5FDcd59ik5uQ2qFk
651H67UM8zwauJKbYOJ+vCYp+NXN8kM8RYYSABlHtDnDvIwz63jSFhHGoFqALHs8fZdMwXWjAbWh
UFCyh48yy+YLcM4RswiwIlZTgqCIi+Lgxo/74kgEMsdE5aDYPrv/7bsU97guGxhBd40zFQC4AKce
gGZ9XQ3YSC5l5tuEMPE8Ut/0vatGP1MVvrDqwR+Z6berXz8+b1Xljq9htde2gsnshGMXmxSCwZna
2A5P5SD64RE7E8tSKdmhmUam6vHd0py4nuKaxflNtR9clbQJIO2o94Zixyk6vc1MZCkl8ycBZ9vt
JnAt0psASEiXbid6Ms1Iv8m1AvXxGxNg1WPDFpyCDCBpO0B+K1JjSxUB64bIrdohMTO0fbKh6ln+
8kGM0kGCGGkQE4e3P8R9dUwqX8zOdhLayEPyl4sGfl/zmJfL5IpUuyC3OQiKB14rv7JQMLUZkw7A
H8UW8k4mQgd3FwxtTuQe8wQct7EOrc+8FpUo3HXYTQGtBv11daBhY22ra4qb3Q1UpdHl2WxcH04p
dLg49lgIPf21UNzZQ2F8pPMyvVrWmqAZt0ZQqKVOA28m9fdHWDZFRoGKnQTinGi6bRbTRtD5NV/G
1g7cf0HLjGTrON0K57mNmXvYaaVFyDzfArhmFiFVAJGSuMrk0tmkJLW7+bf//Jb1Ds1c5V6roDgn
u5yByrztrYWzIyOYYR7CiOSIM/lo5T3TXkYTtVgVQA7quGh6Y/wuYrNlsuUmxhnVaIDjJeUT5nUl
vPd1HzCcn5I7xCYtGf/tNNjTB963QNePHYS2Hvi8mtHMtUiARsHOVbhKQs/Lycs83bFZBpr49zhs
OQTqxx66OhQ4s9wTI5mTwmN9JFbFeeox1Vs2PsxLjYSBuNKPgA2UWxyu9NvkzX5bGvOocruS6lFi
UOeEtGm8VDbVbtNl34lpBRwCK+QXFErTwzCOcZPi2TT4O9dsIsFzE2tvHwIcUDRgjv83jCvfnh7m
/TV6iORtC5LrESLxq2gDTcEaL9y2LH7OFSeHioZQAtPNT/3cW97MeG+6Bt2X5L/BpY04lE4+1ceh
fJHQQGyr7nIwtdzUz7jcdb4KcYoZ+oEpzua1USRcKlUNRBoQbnlr/L6sxqTuUQhzwAdZQWeFg3Ee
5SOWUooNqyGvs5Ri1WizoCOiCPX+nZYrndXu8dfOkkVl/ySmnoLVxIHFXTBYjRgiLLxB03hTirCK
MSim2RFu29bfpWVO7jh5DFzY06wJCeDK+7gbpVkK99BDl191M+Vwxck9i3sYIeRaIuvz1k4lipnv
mKYFW/2hJeNcH8NV7RMb2BhHS72ZsSxzG/uMI0CcGMsKocr9VAEgiL3+yrl6N5Rhw3ElPWRyTtv3
sYiBJkiirjEnoFBVM1Xw9FrojHgf9EszgPVHfIe96/nJNvF5FpMeThd6R7/Cp845htOXKjbG3v7I
sXuz+rSelMJYYoNM2+DKZSbU5QQ9wIHhu25i85TZ4XLK74u7aWmDnIO5DQTt/2W4sRtFU8p1f+oR
0nAQLARTDUIwEyD5J+ltkfb0VSYbESoX/h2y+ObNi6W6xCkltlh+72o0D5moPlH1ZkgDyVM31KO2
33gyMi5dzLF5X3tBm77WCJOTpslllFg2Fy6cK1zLk74FXTrq1zFKCWwRGpuc5iEWnJzhC29m1pQN
3IlOJ8M8nC3R4P6qyAmxfuSU0jWGIWQnh5o9IBisHRPtZWbJaTw1T/dB+SQX+EsuuRjXivJ0i9Hy
sPPmjBJGO9W6KrWcvlaLd56gwRu2rwi/WtMX+fM0wOMzcSqg89OWCUPTzvq8PDQbsRtjL6HShyFd
B7LNDMj4dN/UTj52H0iMFycFkdWglWn8WiD2GZGMRlSvClYN8k1giiJUrbhz4+0qU+hgsr06Vsto
Kq/Edcm9Njz8v5qQlL+jCnbIuvuy4pUyuXfXYiNfKRDPRtSjALkRqCAzr1k3pw561wtfsL3d8VAV
E4Z1VkT9KcXutg7/BzUHfIhSGMnM5QkLh5vqb6NhnWPFAOKmBlHpRLpd19x4Ji0V1IMCe8mZK5RP
YPMx/J/oH+SO/4dUmAA8cxEBGZNAucSDMJlC2eXyCRytHfJ+bq0eij1OfwTh4vtAemxpKHoWaDKa
f+tj0ugsH7nQq7HFIkELmD+AIQELjc4oM0+kcC3GHIlVbyqp+06+czcwr7h3w6/r7VBXP+eXs5ly
FumdfX46wH/QDTK7hyXjm2sME1tF9m+FUBIjKTnCuTocTxbprCDiQj898J1WWH0OIRB9/YQMxPt2
akI8DnII3R7sEjABdSJ12TG6Fw9TMCdg6Yc/ko0I35JiJKnNdnDDdmjXTAfQ0CIap7v7KM6sb1/q
zRktt2qSDvhiRhQK/BAJUlTEsnMrt0Y7rcxD8QzXoa505kgmBCdV81BOqW4vycYyNn9XcpkaUnIq
az0dKoi50yw9swTUpYn2G4vCOzhOxTER32lR3epkp+N1fNzFwZNS6+LA5nOowS81K+Kg/XKEuIvF
/ZQP1Q8QcvLkdDGWbCdCQ3YpvhdJtpjmqG+kAFJ8EHwr8c/E1bKbOTKcago/H7Mq/gXq1Ba4Q+kA
VETTIq+pLmMIVWpFY5rFSkYfm0NqlAzq2AlyA1nBJYrT7o8iQzzOoWURnRjzs1meJXlz32S+rbZZ
JgFxPtuwPABfMEEQvZz0SaCbyGft6w/8haaYL/sFuVXCozUtY3MzHij93QBJD5gZVokhsuUTqr9/
zxrZz8oRcYojE8Y05BwOwQL5yLW6e6mwlt4zT37Mw7WVL4GJXwhDgHgQBHwFtjBhZDvXVD9UKiax
Qzbqhn3gJ9EJOJ1xVY9h1IFRzBvybrc2YxO23D7P4A+P0d3Wnu7on68iK1xqRzDuU6/pL7UbCq1+
3vlE744CGXDshBu7vqrIMLYInYk+xCOJb4tgbV1aADYU75YiNbts8b4P5MttX2W9+N3N9j+tBIEV
zOp9lVT3hLe9Rjh4xiZCFDCdxXJjhrhec18jwdm/IPJ2iMcm8Jves3Abozt7ourX+9TWsOj9s2FV
pYEPZQpXXYfCz9JlkR0viA7OibNVB8LzNsipGPBglpAQXJAazy93sYTzL44pe2XNJJExt0x5L9nm
rC4Ci1Smq5rMh1vAJyyFIlYsubBvtRkU4Kkpp7hJBe8j+tkzVdxif/sQjyTU0vXXbZux2+vhscaw
gMQr5zAx1IEusRy/piMImXSnoR0fegxTPGD7vD1ShCbSQT7RdJWGMkuIczTEo9/msCEEAhUhi9An
rX+vrK4q8R3/TZ5yNZRJyahpNWC2M0BU8k1FRf1L8FBZZc9g/nNEE+JuhX2rTQi1Ez5MD/heQ9kC
uV+2jvF/xP4pBPAj+V0bEnEhTsV6zOam+gZMS/+kDNVaU4RGFBeEzB3eSQyKRDAej9KpYFTvRJFJ
jvzYjBuTFc0yGV/z9Wz5KxhaoHFBRD6FlHL5LHyiqbmq8e/FT0wLBh4FRQeIE8peKmdhwtoLLSB0
vG6qO6vK800qX1ZDHIGt11Lcw2L9/b4u9ep3AueVoAw7vfcWjA+AVoWtR7aKWXCPSyrJdNWesBaC
Fw96xcWKHAyxzXmPdXhn+vY+40VBmYfYAPQkrMtFqe+h0N4Rzn6ow3elQcHy0B+VEHpXlWDh6RZm
MwpPjlaq3t65ixgPKVyOEA5QhmyI3ehhUac3DUQZSN6yvn3we35Yo5AxDiYJgg6aowf3ZIWb7d5P
c4sgD47fKBlf6BZll4uKyFPKfWtpcvprSt8rL1xOaeIv3W4tJZJ101GVs6M2mIPCDibKlqlHLpi/
Z8g3B9m5oPLBtGCUcc+tq0Sz0G5MN5TTJpeIvDRx1jnP12YEEvleS29AQJkIL0VDlbYu6L4KaAQo
zTguuccFUoV/vS/u7Osyog4jZsHhG5WKhF+aEBvqsRYKdvvcMhN7eoqOrIcUESCzgV/Fn5RyPNEJ
3qkpLzRK2eh4wJXKHRn80qKleufJOF30ZtxOjINJE6bmQ98RzB0264cbbSgyXCNTlyfqqGkqbHda
82q20nDBHkwlQLf1QWObZ5q13nBg9Xm1RVxb5kuGDn7pqDS07fEnibUwz4xxTA318KVEO1KnzxbM
uZKNbZAK1GZQ4Sm05gs+JdyMCurVgTJNN7X7fSPZ82miNPk/Yml2f1xV91G98AfMVzNformBW+xd
H1Cgif5ErlR/WzPXtk/4rlJoUhbFCTAX7xUbH+HeChef92SDl927uVnL568u9UWMMNyS09cYhiXi
emZo4+kFFPfOTfb2iktqG1h/VYq7HcLczXkwmMdm22U1aHIjD768xvVqwsUj15yX9NztLMaNA0HU
ASmWa5TM+B9DfVZxS4xwP+7BJu1+zmbyaX1ipQBwsz4WPUxZePZek+cqQbN2XA7Tjg7y04Gy6rbJ
FaHGhMv15WTLPe+sbzJ4ec8bvI9dMVwlCvTQ9nuVC538myK2ZO+RrH9jJy5ma4ZqWGHeOgmp7enx
Yl7rwTpQjX6Zh3H7sPXWwLue6O7PA3zyrpiCEzGWLHXUXcr3Jk4G8p05+XsjIqyG9EdpGjSRjQlU
8B39q0HhVvWVkUrazXd8nk+q30yqSFqFewptFrbpFkaN7DSJjSy10BhVQGyc3I9g9Li9Ea1pnQaC
A1vcKL86rrmxOEqPd6fzuD6i+TFb+3GCyl3r5c71PVIaLz3bWT76rz4F5oZqSnggCV2gkXImJICi
k8Dy2+1gpdNlwncLwU7u3SpZ4q58uq3+3DBZxVw1yW8yzlv7umo51dz2/TO6dycGY/LHcyA43gIi
LwhEvLvKIuop9XyIibhqCuNL5dv618ia+agllKC9pF2xbHFrJGKYPSD+hR6qzf1zJ6wb9KYAsELA
czGn/D/+khNpBxSNiT0dixpAyugVnOUcqtincWsHVB8LUkjkGCoQemPnCNpQFFj3BR8YM+uroOBg
uUeRHGRvVGl4gy37v08wWgImRQXK123Y5D0T5kHRgfn/nTcmw7RHpWgG8Y7PZI8BlUC9jmlCc4sr
bgc+XNi9e8RaTK6GBO6mo5maMMXDPQqMAknUiJfOgcczpQ+iVv34tqjOXw19lf17GRgMpfOIrR7P
MpcfCeG8pYXFQRCzkZY+K6t8seXl9xKJmNuaf5aNgYgJpy4p+PSvyXU2TYU+7DyiYuYHMzZShC8a
n3hVag/QEb6VwKaKjrQTQZXmv0CGEdyN3AB/aZY2vb5Ijs56Z59cBE7D3Q3cMrF+npQF6EXXHd5w
KT2K0iapxVYmL0Vui8T2Z5ikRhTpDScX4fS5PnWQXj08qKqs6smr59iK0N1o0lsfb6ExhqEAUIyj
uThJduSnsSIx2w7dUju3TqwqfcmZQazDhu/Nw5JjOOEf//H5HwdqZkXT0EdxzlxlW0+ndC1fKzcq
x2ZKSC8uxMjtVkguBHUHNSmVEyh6M+jVdtTPGWyS+oP+v31p0gnQUAu/GHbLrg9moZ4+noPiSxDF
PWLAbl6sm0VDltIpyAL+iG78GhEAcCYBXk/Y2MnAtsQbP41iDLkfZsQlUSpxTkabCjXoZAxV3iCB
dFA5efbBDj98l3npC+hoPmgHvIjCXOWfbtiY+TRcVjYGZI0Kc1HkGPKvJ6gqTO8KzLlE1bKIUQbT
pp8IPG/+6Irvi53WG6P6FxpA5FoZPbqwhP8LOQiCIw1JJ3BRl8JQMZIpr9su7XvvYG3IOkIniQ14
RECTPxb+4Gg+K7hd2RMTg+BXzCHZGthQtWohLrUG4KccLH/BThHd0BAXnCiK3cnVASHGP7plZpWY
SfNqxI49dt7KmD+mfj8gNzZsi+bHUntdyGzB9nk9+Iw2JwOjr5XBbJvCDCwkYwVKHoRTRIwOF1og
z1GQG5YVvRE3lOnFM/g2n47TN+eJTbSQIMgSABp3Ntob8GoFTTTvCwpgLfZE5QzS0w9tepL7YlgF
YZS6R32VW+hb5+uKy6+crKa5FUJ0CsVWgjEUnK0QYaYd4nxzeAthC/ZY3wVbEPNB0BqPGNWP5sWi
/6z6BBtPdOGnt/2SXcagwPiww05helCZK9zS59ixkMa5ugogsonD3dUuHd+ncfnHt0EEPbSlVqGs
esvA2SWK0CJtivA2qn5rgfbiNfchRPzhc+Q2YdSum4uIJb+vGtITniY+oj3niCTeLxKypD39ffzf
lgxenuD7NnQ2pZYygklka0TR6e4lmMJJXNoIXieRYlWqUR4X7L5x4g5E13IAcC8t/GspX2pUiOxh
W3H3G64bJxkPlIyLR272xi2419Qvn90A2JI0xGC40kNoIi4sOjIghXrM6rZKAzoG7Iqh9TY/XsQc
cHU55txaOJCksyXibqkTntwtA6/iQnjZzyV5BEk3a8yKsVCUaG0ZUziZx+c/u6f6xqtpprlBWeNJ
WXNXqMnH14zIZjsqH0ZVfUmHYHEkE7Cl3SXFu89IEiCeIuPNa4sli6AlLM8JrxyyPiowAm9ZGjdg
R+l3aYtQ38YWjnQLakD/CGMjcP+YUvRyhssM+U364TZU0K8T4ZZKuWSeoBAPpKR9I4snlkZoejz6
PsQ4uO3dAmHCG0bMgjrpKZOytAr8V22rbw03DdI5eyq5R7pz7bj1H6zI8OwpKKhXaF385H1tkBS8
jJfkzPzl5SWwZIX7dzYuthVzF8aDQcwEJ6vFSo4122v8OqULCm/mtHwTyZ1+kqhilfIPcHhh0bKd
GWwmS4ZfdKQifrQSx9mXTLIMpEumvw69IfYBRaAr9fkrWC6x4meSyvTFCnGPMP7Jdw5YIzBtiMXd
yW2cNkY3ufy5F6E+jfOWNwuGDrslwOo2/Wj2i9O6zdYELQsC+cSQSanDWmO2KdD+UJqecnb70dlf
kRKMQYOMDQ7y4zG58qbM400ac0bHVfn4q7ogEgGp9JgUnpnVC+WiAcms+nQHla7GgXytJqfOL+iF
rJ/shZUvB17B1p397/GUd3AuOeTNicRz5U1MRFf18GHcCUYop7HJ5D19eaMg7W/Vv8DxZa7OlBWC
0juUOpfMqig2nqkwuOYY91bHzsPdn9UE8JE5NBbb40cKaq7gGYpenelkuTIzrGd+0iO3vLaWN/wz
sjiuZTxCWkQzmJRVthnYzrwuj6ZKBd56pUTVsb2aFBJ63Gc79AeSfPlb+6nK4e6THGmNOntnvwA2
xZTWysLdZpFfybMoPhhksVweWuLZ++6qjGz4C6mEyUJM1cSTrotX5Zp6DXDN6QWzhsBuKrQ2EOzJ
iiRi/DYWgbmBtcXURrWkiXVYECP6vK04IJPiBBytyVWiBcFwQkwG4W9hPr0sc02CRTvdrfk2ByFa
i1vx+J70WhDmJtt8r2Zvg9MJ+yW9qSG7vA8quwXF3RPfHuFR8knCVf0tpbTiPiz0gOlX1iRWv2eI
2B6jfozX67k/v3P2pp5ENuG2a0dLzTUH9QBCGhAUccaJKfuyS9xrkKI2OSreHCYYpT8ljsXijQg1
4nuCRyHLZu7dbQK7ff4fZadkwbDcHLcMNGczTxBi1Xt93bqFk85ULrQh0li87Wcp+BfHunbGWlh2
5AsdCnAbMT7RD3O5w3SMUN7GAfIfTZ6zz9cD0aGHbmxUz6NWorDG3E0SjjBfvpwXt/yrdbD081WP
xZKGyxuU8FGz5D4ED9/VDN9Ooj+yzBVDRfxFQO4lXrkcj186ErjDrA1gwIg6RQQYYhz9yEKVazdC
U4E1zj320U5MfjeS3YvTfRAgl/UOa9V4rNnVrELU6UOtWtM6XKR7jpS9N6gG0j6Jp59bTX7lVnOe
OqrXoVBkYr9g4OjfJXPzJCr0g5J5yLQyrQpxbaFCsQ0MQSzXNBTKwwQTB0ZPd0cYa46IBTIE66u/
2+ts9Ih6VNAI1mbMGVq8DRfazYUZ6d6e2icmXNhUNoan9cttRsAKp4qktjMdXzlZTJpGVlZ6v487
rxedHV6DBoygRU1cCoRv80WUIsbA/G+4MGOKrXMk71/VcHPrlQvZN7FdgfyXR7wdY64HuKMcDF4g
hjrq4WNVPhjjEvWBgF4jASTDN6fa419jsrp7WhZSzLlQYW+iZzqZsSjy65pnNqgXMe1Qt/0AD1aU
P8kYgmuGkLODFhZGnCryU0FVyQc1+gIKMmx42IgeWtDUC3FvlDsmLus6Lxwp61hcOqn9dCw4MMoV
+P8BrHEW/pYN8Cv5JOROomQIg4IcSLSKVSyCd1h+ZkHLaPo+6t2PJ1UBZ9LBMPs/z5bfk3+p2O4j
Z0CIT0k8ehsaG7gV9EArbUOmyVowajJrDVCSg0taXVmnBbKw3zGGwixwUxFOLuctXMf0afg9hGkm
q9D9O++CYUEpUVDLL5Rl1kkJoy27Ug4kMixGXdirxdEha/DUTlhbMQUoEmNE+BN+C9D6sMnPwqUu
/YlpH8OhiuvjFrFFx4v7CBvrsM7xtPQulu65lZ5UF9gFSsclM4Eqj5lZmoawG8n/s02UmUNyXydf
ipgYT9wX01NU/4TqITHFyFeC2ovU6dePnT8xHgHD1FPYUQiY5FndL/JCcSMqAUpf9jTTFSIQXqvu
XSOCY1QQqcv/xYX4e3RFgRmyO0Wn0ku91C1asT31/a0Ap2XlnjUH6wGR00JFE6OgH2946Sute+il
j7eS/XdIytmf3qxquezPe2DoLJTI3CXEFIqVQWHV+x2aDpUfo2wtII8IrjimaUDAhBulYrNNJOtb
4s1cWBdvcuGwL+zAsE1hfmgpoDZ2V2DY8m1Vzf/pI0CjUUP0TLiEVSLjbSA35LHC1O3kRgUK0zdc
Ly84RrT8Yo2AiSGw5vt4CkfFNN1P5Pfvl9n1dKQmQDNALBBK4hASetnGqVX/pDFA/pN5UyOVmUYE
pgRJMpQjhOqWE/Xhg76Eh6wAYq+E3OjSmFrHBzw/MugxgaAOHm5SqD7il+8HJie0H5tzxwJeJGfV
N8o6Fx6QVGsi4tH5oNxl0HLkM9Gr8FBFnK7fD+ksnHFkRJBKRDueWr9tIm6Pg5AJqgXGDDXWAzMw
bdMaZKlyrbzEuzO/5qfjtjtSnVSv3RI9cQ4qJGomr8px7rCUCQroBp7gScTAt6yn3Abj0MNXBIwQ
fduWkhGWeyp7Y5sS6/uuJvMbbZt9NDE2agLzmg9ub22EScizIWQ8jx6bGeRqIOweVJ67DvVCKoG4
d+/DIkoVZuanqQZZvmdGnYppisXh1bhGC+l4PTjFXIuMevIVSjerMNBpDzNJWtC+GEGomR/2KcgQ
XDlNXtau2xVXx+x000NlSdIzXeEElni8Whxs2LluuMtyw4i3AcCCvoKFPJ4BHWVuUsmlwz/1Fd7X
R3dXJGkltNp9JHPjq8YnVqF+1vNxjd6lAZ9qqtLNNslDfrobEbUz9H3s2wMxFI5w5NFxp3xrs4gw
NX4AA5rz2O46q/lGLA60r+JrLWEjqEd73LO7tzE7IGvCiDCCCvrw0rrdtcFe+sYI82OJn8qbshZw
JMBC5EoziOiz/p7z+FMF9MoPFn7/7A+ZY2svMVxLB4m1PVEG8eio7yDvZTCKlhlJVGHy1KU1ZlUU
X7MW8/8bVHBPjPYzV1UDP4qT3DcdyOjkladXb8kGE5he7V6gxry9WDsjGhVmeYcJhSBer9M/oCnk
84eA6jh1V50ioTlEvGcgkwWOIt7yS7mx1JockR4EbWxVi5oFJ8CavZr1ZITZVFl0lHeBEztf075s
IlJMuwVWBhVO9WOSkP3jG9n4lqzRiRswPQWLsL04otLoTSHoXKjny23Wz/jQmNikKlbrAeCD0T49
nmLCa67tgmqBxpufYnZZrUefFo3gaepOyKW6pqyKcdiGn/L4tAYh358nvBzEtSlnCnl6WYubN4dO
AJUniHEnIn5hwHPKu/TMmuVe/4rT7YGqLiotNv23V6UrBkfUBe46bgeQFDgKR5Z2Ms625JVYArI0
wm2eUnmVemCc+rFPCHcHcjSvlNZHgcRIK1XfbJvFRtW9g16snLM6UAL9jdb65ZIov9TBqiPWcj+x
5VpIfQjpBAaykxz57TliHsZpDLf51YpHbtMZMC3r9b4vTpVkiarrPiMuKXvPcc2aSnF+ZcSp264O
iQAPWAwcfrYQVzcFqQycONex+hiBbUsRWgs746aNxTg8n7/2eVc4TeTsx7M/aWT5UyyrjgHYcBz0
7pbYgc6F2aXFaR6AnZVrYi4KunsvvzMOegfbDM3Sm8K6Sy1TOUfsoiud7aKjbeTwU1XJCBKSrWzp
mjo7Hud44BjkX7r3VxghbqAqF75egYKXCrRC9DwkaDe2nESBCezd5zANN+FzHHwNR0qItt0k7mmB
NAq3wglfWaw/+OlArLUG5OlaK5fN8Lykl8xUXvOhsphMzDi5xL+HYO3+mcp++kBD1UCTIzkwRdms
oHlP8dHdHmZTX6P9micVJiGks3BVdQYpAtbIpBdelHXzsTxvpNStdFiSYikXzFOTND6ghZZDaShS
SPZZgSP/XYeTc+MIK3ZLALDqhwjliicsIKjkUb1B2M6wybtR8RlAkygYtMlymjfU3RkK60PSC8DG
S482byFOpJFc1wpRrJc+muS85PzgKigxkJoKawjJyFwx9GjFbO8rBaDJnx9NUK2SKt+JElB6tmFT
gTEjE+GZdjSSfWXhFbLRYOdFtOrNaoANL7PwUDHYenS6sWcTF+yDHIU7RRvJ3bXb3Gt5lRYgBm5h
Vgfs/u9CCdb0tNdNciMcpW2gHa/pdX/BKq+55E8YaiAmt45T3kf0KT9RfH4PKYHu1Ch8IXSOM+pj
krKr5biI6jiSkxM08y5l6iqp9lGzeC2RTGBasYHMfuO2GEvue9vVlE5g7WehOE13q3SmwsAvQwpf
6AP/14NrYEySgpqyLJxfWnY42v0YiIlZoxdRX/6XocUZnov7jx8RaYG87DSc2Fn16H+G0FjCrXfJ
Wx8oyc/k8S8c57U2k1HUZLUdFHwEa1ByhYx68wWY3TSLzQpzif0oHcVY6f/YKK+x0Qwwl+biKNkJ
K5afUnHoDiKSi+2U3I8ohC1jLvXY4sdPfXEQXOJJ7iEDytWsylKite0WfTJt8/0vLFa+IqSCPLd1
vsmDUSoP2wF2jYZ0FdIG55aKCisgpvC4sM61kHU07wWzlq91kfOgURhTtUUe/IOmPoWxP3t+7nbl
xY6uInISWE97/0FtlPwouSFvaRYsOLfu2/wYntgo11Pp22Vjrent4FQb5oKDdPObwKNro8d6i3dW
RqDnbkYDZCcQxD/L/Q9kETVuRyGOFKF+1RZ8iWvRM0Hf4bbKiqm1NTpoysd1qkrm7I/brxRKQ8z7
5yAp9yUbVwrAPxgqsGyT3XdfpYbiQeQhccjZITa8Wtyg6S67HbiLYNeZhESjV3+JXgzQY01Kp/UN
okoRDI5gPZ/3eoUnqUV+yakmNCZic7q2etkEwrRH5QjnWiYiSsSZyPqv/oXOhG33/mlglEW8kdKT
PY3NH+lS4Yjb8gKiSEf0DIbJnZD+nkchkBaVlVF9rfK0ncHugTLJPehxO+qJpqlSf0V4jldRWGzT
RhJj4RViZDxjV55MsETQ115+PQUP1dboYsPe3xAPcbfLoO3b3YdvqRrLLBU6JFFzvH9cS21MOKfp
iuZLOCjXKOa37/yomwX2BFT4Sk5e7gKv4+3TQnbCsHsisMgm5vLm9WAqXxRAxvaamMcZEMarAX3r
obx2J8jlEygbtLAGc4G1MRX97t3hsI9To154rm0+e3QmsZ+31jgsWX08/EBwKNGu/NgqP+vQHhYf
cffuJSZoTmNq9OscV3r8RSrpfKmCw3kvXikIGy5cVFESl2O1sJKzvCRtAn+wKBW/tniotYRVmXTU
8dkPp9J24EwERMzGr2j/pbjPLeRTGYmg/0Uaj8hnyDTYGCuUHtqdhUJo63GfKnLUvvBJ9xlphyjv
5HqUz+C1RMkkrFBao6ct83y+lm5GVGLmieO9xzIeOg3XTFyHpx2HlXOHMOxvbAi2wn9sB8AaLyVR
OOvGpt1faS7fbDbW9L13WnvPH2/zeMLjaLfuRpvrRwWaSI7cWhyqNtIPVDtF3rxotQfk0tgUgZH+
mSk/IUmscMVRY+fG3jfnG8+HZ6Jeh68aKdnSZja9qPSkdRtNhrPQby5+JidHhe4lP/YtEo0OESgu
wrE9Jz/PdUR/zYQViZbmORaDQ7TDCF4zhVoN/DeBTg34FLMlEjqq6oS1qZUkwIxoLdCUltSaC4h+
9G2A+60QCa8gEsQvZxseDRD3sYVF81Ys7u1dGRhI8TpRU/cMUHd0Sow2iYHD5teGhprlqsuYw8YN
+pWY9XShThwtqv7SXQbZYNmjbh40HnxlA8qOivg5GLv20QQsnyNa7Wi8b67pCFhdYQERfpizjfMY
mulBmPnITheuA9mhOmYTap2HQFZU/EY1GyCBW7jLLZYhTN53ttZKWEjkzUbQ/UYx++srVKwQAgNT
PIFOUUQ7DyxUFWwQxIe3YLHMQbD+aDCwVxkVkoE4kK9zs2o2C0DATNhjCxKRi5rBQkXZiU5fPcL1
Lgo/jlALFnJU6izAgNKU5zZ/ZVmNfXU6qFg0/mNVwCgnIfUzWTTe3UL/zkXhuQC81ZdPDpHBiVoR
IcfnxlJlqa+2NW9eGg8PCqXdoKma2lpnfqb4j98LernVCliSu04kCaJcED1ZdUqR2xxRpDCH4Zwj
BuIyAffjmqpmExVpQWOORZgMidNt0WL5o3wOQ9PEwjBOn7bROqSNBELIXgzpKR5+JvL9L0+TLQj9
i+IP7KaI7lAtzakPu0PZU49U89NW2styNz4FXHCleCr2tIhOB+Llr3CySPb7y5CMX3qRxZx4HZx8
TPMXVMbsvJXYz4wBsap6hB1ADqaRYyi2jW5THfd3s9csRMY+m6anhiki6L4SxlGCPV37mcyJvw+1
Wv+zFdxU2qHeFP4euQ5/+qTkEzmntqEu65s3nDKTWgLriWxhb/lrukni3smgWpeMNA4Y6hHxh4H8
fgqgos0nQAJcpHiV97SZvhG2qKu1pYnv+jFBrZAs2Bi+JPKYkuET/hnq7mI/K8SQ/8GQN0YJ7VAZ
xHUKtDG33dnv5/ObuCqdv5tkaql1ZQ29LL7q8rO6fSUOq+QhhGTOhNhVqpVUE2R6Xpqzen+T5EGO
a4f+D0x9i2gZLUPJC5TQb0ipjjY3rDa6IpiQJugjtcf6w+LXgHUHPiurv0btUeui0ZO0r6VzQLNx
Kd5uU2J55ZdiqRx4UbeKygrx0jnlXH9S3/ccf0JRhY8qgkz1hfB17vUl6+7TLByfC1cUDjLemBzr
YRQ6eGFjHWJQku4GWgMY06rRkmmUSM/Wz1jFyqT3pVc0kUoCKNS+nxLiG+av0ui2A1ru2ncrFjTx
Mmb7L0d9dMDcrNUdTEyfnzpM5pAq3dGbWLiDbubmhBoj6OLCH8wK2KjAoHzp2dmRvLx7RBJMyrCT
CZumg590aTiWJAES5MzkP5CrlydaWlpOPS3kJowiTBsqdaCf9RrgypGk1xfIH7sHX9N/l5MgBRZl
xaRpEibSBrZwR2ufl56YtqhnIdd8+/be7TfGwxmFnqP3UImV1osTpT5fimkA7gxe4RMgxfHsx5pm
IwGpQgz04F8NkBPBjQ3HrjG2y8M3FrL+dPg3SQkWYb4LYUGHQEocxMBg44hG1QEtbVLjOswZmdaG
JI+cOJbHPUgFpbUHQ2XWDIC7p7n267fiyxLIMRqiZvx6UG+ARgtgKz6SFjOBx3DcdhXvy9Zy2Is/
fr7BVp3/Rdp1SM+g4+U8axSXm8HiFAeIL1N0ZBV5ZzBFHntOxvcoRyWgiXaQ0j7k4RdLJEUwGqWp
QDVI9Anr2wzB7MkQPNiKjQtVOE/K/XlXMT2JBVaQl+SHh2bg3AD5aomBDfHVTIjEVsX1QuU+8KwY
CibGc1468XbBXXmHslBaXCqZiQMMPY2sykQCpsbof7Y+hRIglx/TPdBrxRyrRCu+XwIKYhzjGKy8
wf7XLEgaP4dfGnPidbUwUdIh1+GruB+HMxHUa5xQsteTbUf//wTQ8v4W4PSKIyW2HdMCHjHnEOA0
RK+A/lNmVx+elM7C7/R4TAf6GdnCnNqPGjxaLJsKtAqkI2W8KE2mKkNftQJ+i4hNbkckkXK6RTZH
JrFwjW/bLd/4ED303qXLFSyHdnqjh/WAthwxO7kgkp77Usuqr6Kp3sA4GF1v0YjxEV9zGTcrbfsK
dtfIMexSrXGBX/M3k1KmdJ3bARVGFNGKGMeefPf+eLE8OK1Xp5loT45ZimVvHr/TkbtmoCoFl4Ix
jtGZmwqHH/uvwcNiKJld1MUOOWBndVt55w+SEUU6Kw5OYYw5ThJgre7B84IIwxiwEbusJWO4X7dQ
6OD2V/NiujB4dVLJoqYoIeEHNf+1IIB+TYZBwN6+lUsK0LTAU+Xn+eR1AmB+TahFSKhKc94LjmxH
ZeBAaURdo1guGkjEs7A9ljM7x16sXV6/G9gznulk6xp/Uq/9bJYrV8XlZZx77Xj0dau47TU2j/I/
rcSkRSj1JYUU+UfYLcSodTyZsY/2Fsg1rDsjVJFsxNRevfvGnunUbIwReTJK0KhR/tAzdxZ2FAkE
/NWZb2NaMoazk+UZu5VKWYIYIGRDGi6zFRxv1A/Bk67L90hLsaycMYcvWuut5t3cmPF1XxzJq6cS
67ErGeK5SB9JdE070BWM5ETfIWRg0IqVklB1fsBEunOC8rNxJQ3WQXmYIh9T/J60ZP5+wsKyRVRN
XpnWHkLN9kOhwxz7jsJt2h6Nc6ufvsBN9Im9SDuxszDH2bp2LwvtG9VQNSklvwrA/1WJ+aKnMc55
B6LAgjZ9fuut19ioLmnrXz6FaoBjE5eweG4InFQZBx1qudWrd1Ev0b2XrYpnPa3huLuKQNb3+uiy
t/pd1tiAWsv1HnYYpQgNVTUwVXvBbs9qRE5D1fANvRmESOMQzz+e+hZsJByM9N2ExWhUnKJ3dvFy
ESdebS8ftCyGTN/kaEH+6Xf/qg+lo3VK6p7A1sXcCkJ02b6kFGj51o+hvT9iQC16vvmoJKVAORep
Vx3YhcYLYyimjk3l9ZQd/1Vq9izjzXh/CmUKCJVFJ7zAO9CZDURrBtJYbmeGXd6DN6ZDcX0lnsC6
9w/rPMxrYcwVajh1ubLdny5SCE35jgcd51yMVgZBuKXaa6F1WsaAdlV/PVhp9dkmIqUyXp7QMa9G
GyXvzSPgHO/1T6G0fsvG2bBygn/dBg6EjrvyGKrP+hEEozsOs2SEWnIILmgeliIXnFoO8BDj08By
JmNBY/1egBXgM333LOyBvZX0SZFBNafuiILmdDzB4/M7DSHDPrpp3RXAiD2mLIjyasfcQdaVFQI7
mn2iCoOKigUj/KeFWCDyhQGfOqF5aSejdgXl+x61vsR14rsRZ7bHvHo80yJXUK0Tm5dL2TClJGAw
kmfWzR4+8zTh1KeRafpG38vmYRlYHgoDXbewopD1/P7hAbDrY4H+ZTAKwvOSbdZXuixMX6vggIn3
fLqo/DHpxqV2zpjg3JaxMuhk/Di78u2V+WsdoSQlmLUmwm6eGE6rfxxif6PZUukdXvkGDHx5IAQE
VSb6HEvyK+pruUnpxhdzsgagA1kIruY80r1FTGZLBYkcHWrWpWCC7JFyYM50nJGr03EM9u+UiOVD
zOE4vdmjxPxsuIYFyoJ03xc6Ok19c28Ff2JIBJC1O9bwUXsgxxvmHa+SjEMJK+PxcM6vhJJ78ZMy
G7I1SSM+VG5U90/QiLlr30HpoHlLn+T7LJLbIhnhKcGjt0wmkRpupSzgbnK17fFTJgeDnCYQsCoH
hU+5oo54VgIllNEvQ2QT/DkiKUz+/MxI7vcZHvOqNKcnr2O7TQHH5scbxslukhUd8/UIO8mBWDvP
cJYACrC13EiAReQV26JEkhc3dRZJBrzob2Bgc+SVvmXelA3toMUP/bue7wQkT9v8ZYuWujgT2FEb
Qh6uLsVJTvEyG3yqEV/d6X2NoOwgnzVL9lXOr35S5HCnDi4FYrP7cW4woflHfefeY0xdYjxvvag5
0nPX3TdFAKgENwYk+Io7PgkYtVqlxa6IomMuR9vUOFX4WtZjGQdeeTniFGmVFaBu09aWlo3OUMUh
ztBQJihCJxPQFCO8FK4mPNf/8n+jrt6/t1A5F6sxT2bKJK2QHg9siSuZ7mgOBeQqiwrDgYcimUh7
wc2srdrFvUWpd9EKExQzDOGgckD8Tm0lz4beZ1ixn6EzWeB/S6zHM+s43ljMpmHRuD8F5vu/sReV
kAA7z4C6a0vph1/TZeP6MGtvHU43YnU92j8Q/gSgEVvs+wFyu8q7fbCsdS7thmoJLkATw4is2e2B
FCpNQe/lIKQmreLXW4BdpAxa5k9Zd5rrh7dhy9FE7fZTi3jyIjFYGZKa/V2c8BBVG9Bx3a0KsM7N
xPDm4vmWSb5Fx7YW+tFsAodb9BTnvH5/cwIqY489d+zf1vOWOs8YxJqjJThAExSy5tY0jKfU0+uL
ECp0UFavMrTxcrjtnMdCenwyDHHv3CB/P/n2/8hre5Hin/2qCb4R++26ZxE8T92ktoBm0u8Fp1+S
lvDyLZfp+NkmaC9wsX33h1h7DRMnD7uLI7dRPBKq003PhqmYTGW7HNNDTGXBdQW+GWnC7vjAFVWG
KpSsHIYWFk8JcAUhXy+4esE41PoeR8zBJ2hbsK0tDqQcPDY8qFe1W4Ea7UqRlUOOKEivox76PRjd
23RexD2qmb+tce+NE8e5UFbvy7SvqZGW72qyIuTqrN2XFcKi+jcTOrn1Je94JY8ai/D8Ml2Ut2Ao
gXFL+SGGLRxTQCDkmDSGB9AxKSBwThHWY9GlyyZoR1aMIyWcBLFUr5R1vz3bJhWvioJmJ38Bz64h
0idPSRTeUiZEDo5KQlM4zKRQnHy+XGmdGKYk8Q4UEmLx7G9joyMzhkOYHTCaaoUrLrrtgCkuHI3U
gJAMvuv++AmGtjVYgVt108FoxYOvtHpdW5vTfUu2pZU1vfcLJTnVUv+cI3Ct8GJLeAazWVoNae2L
r05FkannZHjnQt7Fn8LFF8gezxajRM+pj7Hq0PcMGtPzkJef9pxDgAQGRvQALXFSxbiN4ayF+sT4
cjspW2q1TtV3f+dRlRHVR5jQUth7thfr6E2Ur+gRhhorOEVD9qGvHU9L41V+8u+RdB1SRdbcoiS8
n757qmxAO6cunz5tdEzWo0Ng811NWXwqcNXL3An4Xotkcymlx/PN9YnBNl0cIiOuRy2t0+ta3+yy
MIWyswNPdLceQM4YUNXFdre4B0mqanu6MFcJBlBSEjCbLsyLGEe5PTja6eHF90nEVeW6fYN54qMF
yOyPijlICpD++xyDZKj7EvbFctO4pPE/YAnkFBivnbWRJ77O+ZMuJf650SSun60kVbDjbpf8CY09
EpGgDENxsq6Dy8v11tYGWJkreo+7X1w9d1ahRlsobObIbGfp3jWDXdFqcJXcgrNRuDAQoSFSj4T3
jc40XkoEsJY42CpFAfw8XEkJj1KGtwdkUQ3Qzf/jSWbq7hpW/n3ZDXzUZjSBSpNEnlnzPYATHEih
e36kB9FqNyYZ/TLrRD2h8kZCYvqPgRHTUfHojTPQ69gNi2tBScwaYRtY4EjbWKZaPHE+P9w6spz5
bp5gptD+dv5ZhuWxtCp0O7iLKdiK9S2AoHSwmpSqVdn31Nm7n2AQJdphww8xK6e0ryvncKUEU//D
XNlQwKcWzRMS1ehKJ3OxjK4/+xJaSxkZR/vebx7R49eJRcIFC3j176D3Uc3ZmLgH2ezdxi/Gbcj1
OoFpoO/Fs6FNE9hCdbbCIU1MMODTDnkmBYZkchGZU+EfAF89SjNo1FXkLtboS/3OqSlwrpg0GDia
4Cas/sf0HsEDVPzvFKO5DVUDd4s/FAYGq5hKdEULKdiZWJlQAork96cebo6BiPuJw5art5YBfOpE
t95UGKVyXfXA9zpuuTRn5nL852s8eQE0FWn4Z1WTSy6jdmLpnUeh/x3l4XGJTpwELto5H0X93KOj
MA31mDOSW4h0zNrBYgVNy9k3uA/R606Y+QkkdbO0A01dsBtuf8hQOVIn8Q06QNIYc3WcMh6i1BBP
RhExJk0Q5VtgYXYIovTOh/eV48wFgEFbASodrDGVg2RTM4jZGSgjoGgL5x/vrSLL5qVG50oq3ytu
GlQ73V5m/KtH5mwKpztXakZwPwB5GWEFaubrau3GdLw6efzvRrBstjXyZc/4yNOMAs8VTEm3o04U
J/c2MivHEpsg/c+fB0cBcY1nXAfSbDAk9kBxIkNgO4fq9WdfNAwFqUu91XIn93M1hWd9PitRJ9ny
qKCZumyecMiLGZUx2aiUSrU3NaDzaBT24lHA2KyuecttuvTCwGoVyEKlj2NsobojKU/c8HwSuZVA
9oq8U2xCAxQe6nAJXsuzJpYd66GrJ3YzaB3NlNKs5YxBFb2fAoIx+MNqxuK9sxFpKfDgk/udYwKu
7blL67yi9H5eHVqBT+NeEyS0iYGx3zbLfeCW757RAbGFjBhTnXHaZcP+tdMRrsWZTpMMFK2EdEQ8
Q1fqfRXiPBhdS2ezirX0YnCeQSxPBhbBr7Ta9eDh4izkmeMyEFm6yohgPicFq5lZs9jQ02w/H0hk
9JYm55ZJcRAIOHefHvwIVNOTilPQKOlrvKuu8WqfQokfktRsfnudDs1T7Ohxy/yzex8BtVzMeiUP
Yy6C+5YWAcUKW7U6st60mdu8SZ4KzR0tss5oElY0p0/MmmOIubVLsyIeWA61s2IhetFVs3I7IVNA
QNaxQzSMs/pmhe5c28otJFgHtabq2nWY0zgY9/uPfCoUdZ/UF3f5Lhog/atucfW78eg00qkHJrNF
99mzvZwNSHy61wGeBheraGfBlb7grxJbmggU/mb9v/3Ymm3TkZ83WdpMhT8kKLvVXdc9+MVf0lnL
a3yFGpu0K2/qfgSXUylrLBUmh7qWGjgtIgh3XG5J9nvTaG8LOEslS+w4IPK5Cl6ZWy8fefElDht2
LQF+FdT5CdItuMJTPd8U7Kpj4OBnAYe/zpW7xwBk66KATIMMBvtzHA/IRdEKb9F9tioxC9MxQcpl
kMwWnEVP8mmVkVlM7L70qvxkxyY7JgaRJ+XmHDQlgHwPcVsUJTQvpf+UaPQvq0SPlBiYMniqdxLx
7hF1U0kldvzQqBsgUzxNcO9AmLme9zykgTZ64HGl20WkmgH0aGqEba6NKhs/OlpX5EO36cF6P4Om
J/kfP7fPHnOAhkOQs8XALhAwU8cC8PvNfbREn4ubAKSU7O4f+WPvEhSD3Hnf4cR3ga69JO5rXTb/
+TIk+5MllVYHMd52swgdzlrUWR4tMrVLGAUY2i+JM6mmsv46e24Dk24RwpQEb3Q3s1VUN4822vHk
OC+/P52mjhdXRzjx9Pcl5rTY3DNKM4hPgCXEacu6OOgyAdfiDtoJr8WPMkesv5yzqNV8SB60j1hH
pn9ykZwKSvz9K8JhcF7jMDCb4Mrz0mJ1kCjR7QCjwiBKsgFPnTip4N+SUZ35nevseaErMI+u528S
hMwYxtpjNL/dhJrxnyJgZcNIloVvwvFftEUv+XAWMQviA7eP7HtT302Wc+zPDryWpoFANAyty3ux
i4yYRmH8eoc+nv/Ak/xW2fhjM+scfBdrx3F2iTSRKqbjdgdCJbyojrEf0LmNZzXMSLW1Ui0IeIm/
XcU8hcX3fEy343fjR7a0MTo5joBka1eUc2siR4QSlEGlvNCAWKa3IqTOltvCZzobbJ4P4Pj+6tez
o01Xov8930qNIAkOMPutmEXYZwtfaZ272VDf/C+y4Th3TrrUJsddeplVi6hTLAapFxR8oWN4tz3X
f1C5Vi8biAGkA+KfLRwuxFJxgiTBGuH3X6OwfCDUrf6QtiMnl+UjvQDooJskycPliMC1sl/LPLXQ
jsVvhwdwwDScrivNNhveVkRHBRJcNTyY/xZbz8ulB2w26FMUoz9Ej8fFWN594QIqrO+fZNVM5UBd
xoCeJXpwjiLgC8FZIBlKHiQpw3famezDBQTVHQH7XZRT0kuQQvbDRb7p3By3UI2LjsSCJKLaNr6Z
zYxIEuHYO/fqy1m5Q3ATOpiQwh0XZqsFZcLGXhjbkAoJsgEWKbsinb1ELF9o/HZn2+2Mx35F2lQG
upS2B3oqakjs3gXu1NWlWVFlx9roEGDvirv/ugpkvtMv1kXi5roonno23oIuUMWdecoYHbfZs9hE
x2ZicUUwBYbaipjahNZZPM/KZ0SfA5Ft6P9OOgMGxSkTAYiSvfJccXRLeEFGJftYyRC0KmddwP3v
oLiF6q3rEn1DcBOzgQYa1VRDIjI5FI1JEUIPStOuczB/Mh1IE/2Ajgek/Yu0tItYJA1DmyNL9dcM
0ekFxFBYtSGDyJRMoVtBMAJGCUySCi9KokdnwQw1XsJdzuczlmZn3gGJoEBccMlIsi3ZohBjZySB
uzcPMLDTsG236uRPCbmLDFQp/vvEaUkXGGeU721a0dyqQsQujWStyptKNSBZkichomXxzk3E3W5i
GcaPV3eL478qOm5jYuHNBaf5mbV0MsUCvhoWGHNCljuN1GBZpy3RHmrdZ/vmFxhI/W+Zu6gM1Bdx
CbAqjQTOODCllY2wSoQ20eoNAqG1FtnxUCNahMD4NkXwdYO88a8YjKpWoF/0oZLzdkQG3MvxrpPN
j+v7Pzfqj78nbtCI25uLWh+SBBcVXTbAzdSjJSI6kCObqbdV65DjtsEh/eJxG4P80RX18OvJvHqW
2AkXY0YCArsCTTW/8zpM2WHMriYupZdoc+o3/oHqxqST24HV9sv6PoQ9Ei0JSC3/EM1lcZqC94hU
57t6cE7m3nWrmiJv8yolCpPuKi4QmuLD89RRe1YFQ6htEXawn+y0yE7QRQRp7tcyLzv7s6UINSXb
paR6lpFM1Hj6lTt38s0DVtEIoz9094nRHDhRum/cwft/wdYL9Ff3xnOR+nD/xhCA/eNvQX63SJnz
BCuegmB4n63H9ecbT3oOrYFAlMcrPJBiB5t5GmFJSt2j+OgFrAslPWfi1RORkak2V4yFn4w92H8r
zni31mdUB7vUKZlkN8wH3CDhXkOt1m+dGy9ScNfP8HqcUangrW4HVTYjvmKzfB5LVg73yjha/lK+
n9gKdy/WesW1NTERs3SLlN7WAl8Fv/OaJNo1uMQokc3tOX4QUVzzZhacIUrlgFROLGvkhJNl0ry0
XpuQSGC/Goe7UKKjjRo8048tj618C1h39KCFXEizGJ91V8mExzGQSIbZMroreUpRF3CRt9zsK5da
Pz/i6cgWAZp0jM6DrfOPdAHbycgrxvLL77DBox+jz1dnBIRre1k+Os+62PhPiL4E21EcC9uwBVrE
vKUw/2evxaagQ/uMn9fITF85LbY/5Olp5NPwT5KXiUZ9y+089PC8glT7CrrSOplgI/3CS+Mel1S1
PvvosmRM9ygrsUris/n6CPCK5yAK2vCGxi5VVstsDAgjncvdlUs0s6T2ozo1Vpd30bObhQ5d/nQq
03XlxHSYS5D7qQk5oX0YhMaVJ7jopVo8y368EbIRlOPxEVCQs1KsiQXsGSVRy5/FOrPmardzlYYM
skAwER/A4g66p8sVZGUw3t3QpNcIXaij7rK7XKun+mkx16iyLDgXDLJHH8PyJhb/f+UYUtsWJ9BT
QusCdVbJk5k7kUbGKsacmDA5qeeSlJsP1pOiSDIghtwUKACNHY7/658flkuQLgcCQQvP3mZX2P0h
Y2Y3AwmvTkOAovBhXuhio/W9zG2jqU8gp/fPaG1ktHvWhzApCOnvFgmcOQI8sP0gzvoLPENUIzqn
+UU/eYiBgjaWGsALnqC5L0mELLxBArg5GxccPpevnWXPzZYaGcdL78rJDSBM/+2Yg1i36AfWpnJI
fqT908efGo5El5oAxvkrcPrQ3Fc48xRdJz9tpxh81vKf2ef3mrB7JB5N696Rju9Q1+EUzozXCvRv
bUeDWYimrNWYFSB8frrSgk6qe+Qnm5xtg55xruR7UJmYEVJQR+HGY6SPKmyyi1ogONjM46KmeE64
O/CoFxr3W1V2D10BHN6WTAfRE489q5JDNd9lNXOvcaSm6ObpkLl6YUJsD7z8Fb0XCrIsMFhKBsTX
EvnhaC9DHl89Bc9XASIKf2Qad6HJdrYSuGNKItkrSQ3wrjfODK73caOudOr37DZhf1tjLhEw7RK8
aVnDdnmbHm9Chfgo895NBAdG0TpzuZyP/MoNKyI5HLNCTxEwEjb2CQxhZOABq71t2fDtYGC14fgk
oIqBWlPIp+wuFPuJbnI/yjZvOiCFguI2u27eJEwqziygj/IegSiHux+Qk18MHbi7XKwbUxkIXPAm
HURQXVH9h9JEfEQIsYIb5Dqo0ba01IBzYWo0iYAOdT//sVg02wfWH3h6auU6uOGKsvUV+XhljxmN
9QNLrrA9w9Kq4FHNOZH9rEKaJ6yeeJRueX8oMXFLcuqOEelGcpusZFc9zvJrFJ0xAaQKRPupC75i
1oCh3G01R6/CTjfJNOw/91V2FOjarCc7gtc+aVwMW9mk8urmBfKBvkURLPy4Dp1z2QOsLMO6F6Eu
IixL+5rkgLva34At/3HUABtnIkYFJu5EWbnK51dfBl5cL7TBfdD04YnQEIAdWem+XMh7r9d9k1fr
KRZk6oQQXmyAuQCnqLvepuJoTrtQfFzZMRybqMRm032o5C3/Y3DtQhFMd3zoy/9mH+xt8xQ5KBtZ
xaAZljpyijR+bhyR/+u0eGqLl+6uRhC1ezYniwgaLi6plyRcrnMJ/KNv7bGNJIGYTt4uqxBkKbAX
IUz94aRipBIUbvQFMBiHcAkFeMkr2A4Hk9jx/BQ5rqSTV09ayZO/FCRxPTwOiDWG9KpChPGN+Y3C
qVUojDptv4/dHb55pCl0WkfnH71yUbRLbu5DxgSyNlnxt4G72vXNIuFHh0NTWhX3nXT8QIS87EWA
Ree53p9Pz5T8v32TPeM7iyJV13N1X6HaUf7CMQArJcW6j2GdD266uKGxgSojLOlA6T+YbHIt+gKt
5CvGUvGEJbdbHul0EnMgWr81kyCcoora6QqOVS/2JAnFvD+mmtqbfXAnFALWDjA7OTzpqlGX5EQ+
KWUPszGylFwCBCUaVCl5WItnw3ziKXisrY3TYKJkcIaYK7I9doQzput03l+TzrTd7jt3ggkU1Npl
KnF+53YGhBQI2rPiLLCJF1DpXfakz88CWtgYph+xGiQGAnUr341/Xi7l/8RczrCxXahKxMMf3xtZ
oDsp9JDL94qlTjVU84f9S7EeVexUteicCGKFCXyOopTYJSz5fKgUHYLxOpc9oECFTKEkVAbM9MlP
tWMwcKRYvEPf+e2AOWZBxjBPiAIcM5fufmtJPtHe4CEeAaytYnsrV/rU+7n3D7Kv78NRRC+lpJkB
IPCefw6Bu7eOYReANZNH6Djcn2tiuLvkKcanZjQplOzdBIgwAign/Oa2glbQr7c7YDlSlI+kG8Gz
c7CuolVoX/tWgQ1gQECy5Ee6CNDKC0CIWMcwiNiP/dgScdsBljB0Lcw2XO37D6hlZR/gPZ9t56UU
TBd9rwGkwKyBwQVELdbCSUYLQn/otw7SRsFZt7jrL+9/pBrc1QNt2viUWAwbyurmR60G8vjy0TOl
Y2D5IOqUgVLmZhXgUdnNMGDUqGanzwhncoJJX0hpt38wmLdmy/vApvLiImaXcuQF1fG19xZD8xos
S7bKqmKEgP1D1nq+3gEaRpfYVvyH4uhG5fRn9dbN9s0V1EyfossvLc2WhDeoEGqRsxzZFrhKYuQF
S6Z1dZlQhc+wiaVY6p6PyuXikgLS97s3ZcwE5tjFe6PjiNAsSfUoIAucHDfWk9/5EGPQ4PLBGb4/
/uSjeU5QvfxFCsjmFb48yprHOLxFyep7Lbssi0EK3rFDwnhrebmB56r47vhcaDGRHM/VJzVUbO8j
Ltj0D3NpPi6yz0STWtFxg/UIDgDh8i4u0aA8L0df42vXxKbcBbbpCps+q2p/kHk90OfpOeVTZffi
Vmqplpl8Ejbhiu2UuAWreLURCDuPw0ygeX+TGl2E+wo94jtLzjDYZlXOvMMQ8FGTF1WTWYUqEL1r
e/sb6r9/agerxdz5238xX7xywvfEHFvZ8nE8sEVcBPsex01T7achUhOcWqubzPQGoIRxkyLwY2oJ
OkgJ424UPzDe7zml7R+LrGlCDq8nmtdkyDofr3Di9rkF9kTKAEMm6ym/FBdaZb7LcLm5iFlTfm0Q
jDRnTjrS+hGhfQLj8rYUKrUeSGPI3zyR6qQ1VDPLOaLFDIqUINJ9fkHLF86Q0fx/c9YK50z1hh1g
BCzeTpqB2K4yWsUWGcVQPjSH08YXFotGx9BT0KAlNZYw5BPYVRk8UzPHdp3wQi5RZ6qfAOxBNEoO
AaK/oXKnCFesRuYAV7usNAakD65GmOdQfNEqTg8eEyvvQnVbZ6xP/soZ4twp2I8+lb731TtXkm+r
Jyq/ePtYluywlkTjJBm5FqA0dXAiPWvpEEHUWM2bSDcHu5qpAHGRlJi6wz74usz8yoQynGfE/MwR
8F5NBWwhuxxB1OhTjXFTCevS0ky+aMHgrnoFU/5yLIURXmDLKQogwTZN3knz9kmynmby7ofBKa02
9MZuMW5r/08iPSTEZ+6wn+hpLeGQivCuqeiIjcFMn7hAWq7gITf3w47xGuh0nRZNvNqbHxQ7pD84
R5ndMt8EXseGp5PYwOy5AZr1HzDuZXO5+VMFcrySejpGBRplSoJa/qXyuHPpFQLN581UL4yniM+L
C7T/XAYC8dRJGXbnlU84l6fspUEWlugOaxf+2MeaX2sVygLTbUM47A4QpXcWjfpvclIIc4NoljHI
xOpdvhPstQOyxuSAGuIbZV1dEEu7D6oJN23DKi/rSMuBr5cT77BHYR2GnEWjyz+yHKjNWoQHwduj
VFbSKvjcl/ymmVL3Jv1e2szigjPAit5xEuSAbwOYQJbse7FhzR4Oo1E0OJk339tUbL3NqLYy//JY
9DBl7D1VjoGOwG+yySAd8jKaiLbHcbGc/uWSkU+FcyI4mJQ8nKRX6EgmE4R1NiY8vZjqyVJ3JBEw
2Ivggt9ILlu51TG0Qn0W/oniR0+8pSiTgrCjCyjyUwxhUcDSHNmK23iGYlatkGqyzLKOL62g4Jrs
5PNyQimuxll+332Zm7W09EPsiABBncLEi0UPCRZVAe6FPb9vIVjwTLrn2kDHFT5ayKF9yKg8X4/m
p0sJ63OjXkAM0Gok5fWhGih1lKU0m5gFJ4QOM7POXzJPahxikGUtQ7Qx9/nJfO+NJ5HonK4POeCI
Py7RtfoPMmOP98UF2dU3FkRwJ9M3QcHIUEcVEHIx46y/qcPC/pwrAc+zeIUTZL+OqhGxTBVZNK9V
FKMMY+k9Bb6Opf4xmSI/w8CKY3GOC5kjBJbPlVFUqyE3ZMVuCaKWCNkIPehS92TOjLYU2KXLel0L
6g1/lJVYz4375AB0Koz5a8t1+D37TjhIKgYln/4Lc2JU7sEEmoQQfqfqfmi3KtLk8+1eTl1pbTL9
oBIWOxluE/zGKk+DzjlaVEGQeIkXJO3ZGzVM39dia4fygg7cxATy33vQ0hMeTOCrlcCnrAB5xVxu
p3JozAf147ap84YzYNvlVd2quR2RKnNGjWKEwxGOVnZfxWgP01TxfIe2zVIZmz/viKUqRYpnDnnB
x444vVZVg5ZVZkcegCcIqVzCq0hcWjwRzGTsi+wd1SwWoZhNXGph/rXZRw8rU8T9pBcBaZ2khH3g
fSvcfNyRoIL8+DwPWogrZW1fMV0DaeVLM+02KuiBT0xPLGvOrdm9FGm3LeJSQmR60w+iKbUsNhfz
c6UDnWavf5VTn5zAk5RKJoTRZfeJC2Agl4WijuNtAwAzdqdIFC5SLn9RL16P0sWJ9Ca7+oLT8kS5
ANTxN3DBH0jEa2XdIpJF7xs+i42h57zO60X3TxYvNGlMEWvfWe99ZJ4JH65Bz3x4KMABjPVdrgf2
Qh09uiZPd5S9HkDm1Usrs8HyHQy97APt9volsdyKE3LnRH2OC2XohsIyrwWhk470yCCmVGorZRWx
6Zy9C0wDzKDRiGwj544cMpznMs4klclEj2rIGvGurBIcdr1SuOlbQ0VAIorhFbPLEsKL0MDMJkuA
u8kvCqzbRRY7WKrbiY/cGdjjb0XKlyhO76X5ZruvYiGxRYK2BjtO9EB8mYrsqc7yY0AH8IdqZ+yN
mv8cO/LI7e5GJEox88XKv1/NHphTf1WNJKTilfwa+28PqF0HW4I6CqCRKZ4iLe1qpnL+d4bJUwBF
h2SbJ0fNE+t6C/QThCFZFHqndqEsJs634qPMchN1PTqibKWB+4s9oIB5FeaT69CJYnbLAffEbZ2B
KEeUC1hjZarJtpa1m9ZWgjQ3v6s398DOWnlyfdY2giILMW0p9IgZHkf1rD/qItuytoNAQPnFUUkK
BGgVkKUvqU6e0qJaun4ghAgHem8sajygJjUG8A4heReSqBzc66RCf1yXFrYBplJWRTKVwTPGE1np
K/PjV0m5UNWd6Cyv3rL1jjS7VAsHiR9ZdyLXuBycSPbUWesFsnazSt2qIqPtzLdt2Cu16rhxQUnZ
bVvxY4UNyqer1ZYR331z+ilpoczWprwBm2uLO01gN+6AXQSyE7Hs/H2ROagf72dk9kj3jB2FqLIv
455mgtPdYJClztGrZ2uV/F3xOLZBVmOTGmze+IEmb4Z0qZHiZQ9BL99yJ7FDO86OVkLVFJ7xKZ5o
2UMO5FJVZo4zsxcU82KJfHHFw9Uda9xV0NJ9k3Wim/yYpqIa/ZH3H1b8xnGsILfMlOEEPhpV6Qwo
I4ZWa6Sp0iON3C5lPDmIx7bS3mEW6wlz2S8RxcKRk7UkkIzAbh3Ce7ot+gGoHVPpZb3ptc/pcyGQ
nDX/nspBlIuDfDdqI3hgKMrvMOdSiO9gvkBc+N/lvEi3GO9PuBZ0cBZIATsUrV3XUVO8+qeLxYcx
ALw8mdBRbNYGOOY7ruMHlcKFWc8DktGRRyzQXcyvMy64dPQkS3WEH8NOaLcklZ6gIQRe06bP5rCw
E+3Fq7eMoMEb6wh2KDDOYwvkbdwTrcHc4yT2zryLMicuR9lux7vwlGiP71IN7tsvnLRDjEJk3M86
VjuGysNJbo+T3BXMZcEVw1RMSZzy+LoeaadH2TjCCmErCJjyVWIRbpN/ELwGdfsa492tM/x44qla
JGZ+7z363auT+TKf/Xm26PAnJWRKEZTTuHpF4Lx0yGFE1e8fgwd/rAzavUF7BsHtIV1tkP2M+IQw
4JLuyPUpvhSYkVK9R/oDHjEt92BgkX6q/tDZ91Y5L6haS+a8rjWLE335Y9KNiZXmBgDc5RXTH2PJ
9VDtJHk4RP5GxFirLuFEF9LQksY7TteYLTOCU61DcQsvLtWhZfgb9kH5D2tQPBfr6dG/aTz7Moui
bMOhATDM+oJQ9Rs/N5IfDHsCZiy5z9CKgGwKj1sOz3Y/FlR3it5jffv6ktB4ynce35tWEtbBPmfs
H9WX9HeYuYhCug4KDDlMhA+4TxpxITgZoVHCcSZke9Q64Kvg0tuqcBYRUxa8uSS66FxAioD5cumX
WVobRhSfretWcOY7wNWvP7WgdlKoWBR2habLaiwmqkunZPVkH2B6H7sg5eo626pM6C19nCmAuuwS
QyIMSib8ntFYfT2V47cGhaJqGntRMgH9sxrEuvTBQHGt7bKQJ7b88Lz70KkgsSnf8jT6PqNnKkGS
p4MFicGFFSNoEJMsZKAcknOzH1oGL6paCCLFEltRMEyJ/buk69ZtDe09+TdbFhi2cl1btSVKYAL9
nOrdsCHvOF5iBzwXTDW308GPVyLWTO6jzdTfFr4lF2gKiksSVwnH92Cej6oMpxpR3yHEoHve5vHF
iywnB4uREdA35O0zcx97W7NCWG/pPsQ9X9oUCzkDIwDWzXG7LQhSIH28s2QbB9L+nGT3E69FFbVR
jLaqgi+Knn24nSDOY3REEqD9NQ6S3WpluQRdRkdLsgJDsXZKyKODOnX1FFnbXDN9PE2xLXeC3nvG
5fzOoEIYapCIJuo5rF8c86CS8c3SML/xdEAYC7kTepf9eVEIcYRCAJlqlxVwjq6BtVmkFPtzQcwy
jaiyXRdXrAFOqcrg0p/DiOUt00ooIq8uKPT1J+YDXeFJ34ecIhO8C0VUopr7sB/cHBvCuj9OSooA
jLaubaBqwAgf1Z3QbxGEDi1hG7Lga9OoH8M1GzC4a8TlavpTZjuAs33s4mQLQv5Uk7bdHgSM1xzj
Glbywk6TsGqpqI4KXi4isiS7F16m24232IzeQjpCzTznlq8FoEgUdoKz+hE/UKBMdG97PapmcBrl
nTlnPK8KZDDX06+xzsU6z821ZoS7gWkGIdzXQNSgnawymIjNozZFhJ7fIHBpDKwAV/h5RULxdlmz
LcYYBma9CwsELVE6dYuWgjfy3p23JZ36z+yVq7HJYz+k57yAUlgbHZ2UKa/BInPE72H1ROLatr9m
HPN+OdM78p/DqBtS9+Byecnt1fqbBfP3HknchyJaaSQDgqWT0KxqPQA0vkhAmoiWZBKN6MbX7OU4
MbhSLO+Pt8Lo+l2bvK1ylXRjPfNbXwSJEBled2aRLVK8gdmMWmvreyEa2jBCu2hUMaYAfUcRYPr4
1hgsslUB91SmzlAjksRVlEFKBdARQnnJO0rcomG9ArfXhRh+byzVeBlZncxV4ou9Y9Wj6QZaue43
UFxG5CNQKMnKXeG8SVk7d2kEUfi2ogP2y9CtYCnRzQCCUBl3Kk/RWCNSXaK/0ImuLLV9acq5Bptb
SSBrCxh+T8aAt7pvzDge65l10+d3q+zAG8wVBXuDMcXWTM5QnHwanUvWSj5w6BUm6nJP+TeLzNu1
241repnsa3AHbl5yz1u0HNRhQKS7MwTuAs3TaQSEyytC8t/xwh8C/oUQugomBEueG3Om2WTnLu+b
yZ3gk4s+lRwiKaj2UnhZ8Ulp5uNrPkGZdoh+ULJzqAcKfLjwgtGOH9POvnNz90RFDnID4GGDa1c/
osOQIJqO6ATbgLDgo4M2lMTCGcDNMWG2pLqxCzKE
`protect end_protected

