`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l74IqG3tdCuSyaO8ir/3VT0HzTwCNpl4UyA2wq3bn+o2c1YbtZnJJmc1AssaAZ3CLwE6j63tghc6
otN9dx78pbtNSc2cmFXE9EDDmuqawk0LNuqyzIzWWtuRliovbs2PqzFQfL8YT6CHR3WTJfNtxd6m
swKAPSQoVgevFPDh51nxZmBQ4NViSz6f4jYeZ0QRC8oGJqwIBH/4HplgnP3Y8xAhg86teYZQx6Bz
EaiIz/VY6EuRjSD6u0/CBG3tAsVBaDYJwdX3sXzz3q1/rn4ksGDpD2GaVA91hK6Ocr+U76LkgUT0
+ocAXrKOYKb0kbZLuiST8yWNSM1TC4yRD/hYKw==
`protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`protect key_block
F0GaBxpYLPuTtyhs4iAYqmgRJSAwilgpiShkUUQhMS6QyYsIshkK0A93CBnpLon4hIlGZK14xrKX
ETKmZEkNe9UvyUj3jz6rVCKK0/efs/2RgUVRDefBA0n8KocwcRoS9D/SGCiwFTWBG/guptUJ02DA
BFx8ooA5ySsw0Iz3qrn25F4Ds0wCR+61etQOBLXYOfzeFR4bz91ur37yI3PZ75hQF5KTnXkODQ7h
x2N3C+KReTIVvHoexzlF7MHvsFpU8wg97Wfew1VD5DrddwN+gpNMACOkkks8pI33eJa+SIFQYh6S
JMmWFltVdfCXlkWjq1LdLHcOnh/NX7Dhq6OphwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
i4jiDxOL484aWBLkeRSNU1oilgFU1VF7fUMrOtXpj1Omc91ChH+Kd17GkFcgBy8s0cU5SGTd/Zg0
u2YmL7e4KA==
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m5RnXv3+J9KH/fnKYz8oT49S++tdyWWpS5t48/fLiv3h8xSgmzh17X8UtjilGyAbJ11VxMGOoFDW
r46GGqjaUvFYjzlmNDAxHdl28r2p23tZjJbJbvrRN0XZz4kA3f79wovX1xoZSROGkj54yIdrAYMY
1wkq6JCw1n+x+/PO0dXs/rjWrOnvvJid7Xua3sAElznsQBwZyzhrpXKSy5/KEJUWR/8bnMzDLTB0
FUlcEbSYiQNsOOpzFuD3G5JcWzlM5PprYW/ITHp9N4SQ9YpcJhSwByxRXYtfbATaWWQurRZHoBfz
4PV+vaeQWXXGdBjfeOGlxe5VJ4cabtga257w5Q==
`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gKVvaCmPooegIgvMI+V1uifJOLtJfhdecnBWBzBBcg41t/M9/NitUGaEDi8X+49GHRKx/iteCX9A
zlqZzqEUuk84DoCSf5OOhfMSWCaxugEVaucimv99QSpgaIAf4sbA2lZXnS3elF53NX35v5N9GJVl
Y7cdxJSAZTgrSoFMEHSwKvRgVL+rIsa+lG/KIEzEu+mLPasL4xL2WnSUhWZTPs/O3jwC79PIr3FX
5QpKCOrk88GqV9sDAf3US9jTmEL76W+dcLXT8c3gu21Dgr1amdnBoO7S9itoeVdmw+PgmQixWIz6
Wy0XdDyGW0usbSi2zy0pO2j9baF3suhlZ44iUQ==
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YxsnWZTKFIX3fUwGxpVPA+7ok3oqIpXnBc3gLRGhT239b2oalywx1wE2utRXOyYJJheNy80tZ6Hn
VCqi8netj5k024bnVyw/6TdMjJiOyPVBiAR1ua5ehLmFqE9GmQQGVGCrTxZuoW2zgOFsV5lzX7uj
d7WjcqYtUJnW8pBT2vo=
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F1AXdKmzT7/Tuc3kxtv/uTs7+XwT+BNervonN+gnd8AsQv+qv9o+6MYT5Plhc3C0ILIFoi4I3lXT
Epst5fHGEsu33t2C+Sde0YUYvz6sUwYYka0Iq8MWqvQ6cg6iSLYgugSVNp4xl595XqqSg80QBTVV
fJ1ZoUi4yrSD4QmX6Qd9WZWPbs9xMvs0ewzFSR35F/wcP2FuE+eOW2QrPkj+QALnycJpdB51IPrF
akJp/8vIXFazZw5n0Sz0yc3KWtE/dQ0iPAusP3VLrib7QEbX74HzIBbTmDH5pbR0XmVYKTHFr+WE
oW6l8KLSfET3cdhsF+TyG4/JLlcMnsAPp0KoEg==
`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pryiB9JFPjIMGw5v5QS4kgDRWaHd8nKwj0yhcBmRQljjDu0kG7KVDM07+eqpUXA/1uR/eKNt4pDe
MzT8KZsUoURdZ7YdslPPYHAUrF8/EUUaWn37vO9Ot0BtTfZvz1ZiGspbi6jchJT1GVTMBNXW261M
1d3Gz9081P02/xoO0dsl/viLcCES+SnCGGNr2LAz1eDq4bEjHhtU4nTEwbvrpWw0RUBZh14zDoCa
CESrTKKeoiGVRzVkqT14omRc20d4BOc9GEqPt1Bj78JIp4e+wogPy91ib9cTCGFXMYAk0bNsXsJk
LW0nGmACFno5Ua5X5Q20BMtJ9xOFcN06CMR+pw==
`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rtjBz4ei9oRpf4OHhpakjuqMkKJTyE6RmDesYp6F0EhKtvlBSR9GY+AFUvtsSKgEZ6k0VOVZgg4m
3jVNYspIERAMKqm+FTso3Hiw0jG87Ul7z/IEIWYTkpIyUcjRva/aQuOh9DvAKzqMUMuvTfpSvakG
fkfDYdq0NaddY3uoEJg=
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pb6xq7Vf99Xl7qiIZ617ffdN9g/8aKCrGY2huBrgvi5iTxf9zmQBxICIXeCCLZ5JwM5At0+ZGYey
ymvnzmaxw0Fmuowmy5hfOImCsn8AvE1fFBTeMYkcHzkuGB2IGWGu544XNjrHCY2syWoFBeKvpOmK
YL0/NcAnc5yrQ88paGjDeZ5VMQxobcHt0c7TzRN7TtXjlzbZC61wa1h/GVue14yB38qGytIt9u5O
968TLhMJ12WdiiCzKNTP5H6KQBQWK0YNcL7DHv3jfvjFpo8OZi5kzWoYcX1/R2uQG5jmObzTt4vo
AzfVTaGDOMTlNrkOJqq+bxJDYaAcKom6Jh20SQ==
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 63936)
`protect data_block
iIjzykddONfcrmohy/CjAYlmOODojWKDuAAwsCYDJPgfeB4EJ4xfxslIJLjOuIm15nKXaKr8j3F2
wYagBmSzmrohM1agQW1wCiRYy3BHWbR3z5CfPWCWEodEcQ6bV78qjtTE2uWuk5XYfBscb078F9/E
y82G+j9cTZA4igtDb1mbxeDb/b/uEOnbd4dab9dg3yTmMSJjlzf9mHmNgDDNbMlXyvk8NuRFjC6v
OWaTeiCnuFcliuM96UMZuJQV24D3j/6hU2+NWf2P3xZgVtLggvx7A2EpnbB0qN/ogTsLlQ5QrCNl
wJ3rFJRRr0p6zakys+hO8VZf+6RhpN1Uz4k0O42bhDccWtNAEMsEhfK/o4txToINjjH3hUkmj7Gw
S0utXRfai9rlnSefFNiU/EfyXdleMXKQeuq0UfyzaScOjfe3XgIrCBaHVbX0IeJ67jcZv1eO+1U+
TKamhW9NlylnHp4EKhy/HpuRufbz7UG8rwkU+AX/rxql2hFDfty+Ofi2Gh6jb4QMXnatFE8OMXOC
jGHCJ695JUNIucTKK7GgB8RBoVtKy3tzlY8U2RWlVfTIPFkWOSJPHPKu4fnb0PEO9JRx37mkXukT
TOuGaxMhDW5nve7IMMx8hfV35K5MOx17Cj+cLQteElxGLlWCuhjo2qNzFrOtT0//AARES0dB244U
JdBxHcZnCNQp2LNQl7bDUzKnJkBVPdmDAPKFdZUxMsAhr9OlpLhoZ8jY5bi+mlQ3zzF9LNA0eSaW
QgDTf4H+WMnrvQ0ddzHb++ImNUw/GQn33Ej1Tf0SOEeShj/rABeE1Uc3zk9Y0rE3DAUgU7DRBjw6
Ym088Zp2zbsNdl8sIhNR9gMn+1J4XtaweQ7ZTcZM0QZLXanEhgmjmKFQ7uUoqdm6pUDCqD+xVDXq
7wwBg7d+5f4rjZIjpl5A8gTErdH5RUAnn3rsXRrsCcIfihZOKlJ2U28/Kct80bnMuJT/Gre3D2Sf
FDiuisbBbeKQGokxgHt1Bn43TmYBA3llABnZElkxrkHWpe592zGm+SG/0TF6WQWykzCMIzqWjhgn
Vy/w7kRoraClIH3yWXcOiIj4SXaogYoWGs+ZP/pY9iQlETwoF3Ff+3oaNyFr8OxEd6KlMoqHOEu+
qVeeEQdMT+thVXN0BT/aDZKs4YQhVce0R1NbVabCNO6bGgM7Ib/03l0K7JbEFZ4PQlWmT3gHILky
QAj4FaaHQ7S4zHREtYckkHtermX8W3ONCfOvlHkXe6/mtdUSblIklJ69EUfdT9wyEFLSQ+bHWByF
pRQJcPYEU2IXOXXyevZxBwd9QBxZNJZbqF+LdEg3rKjWzCAOFFhwkZrO0owh5e4vkZRoQjD6pBn4
DHV9p55Ivm42CRY9PMbybYWlqJuTvuQNO1gEcLwcTBBxq85jHEqq8oj0IO5JIGgFeAniqpN4qtdx
61RM/ZYuzUpx97rHH2WF2wCnr6SJmk//1viZhz1FZlaKk1AuLIrwkbS7R/BJYcgEAU4BYGURxypt
h4SwmztxZ1MFbdPoPqsOvoMQ2ArgPXNfeC/LnMSQVJ3AXXriEHN6BVVM5fGQAjeSvKDrLh/ICayB
LRTph26RxZP6vb+ByRxgx8OwKNgk9g8buudWhK4PzZ/7vsAE8iXvRdmFSV9r0wdaeirynyWjJYhQ
rW94ldbzbsQqQUdcsvZ2+0MFXgtSw8aOQo90lMevSYuXDmKMFOlULaDxo5eoEbjRQ8lHr+7sKK/y
1RIlGKcxz8goBQrUfq6cX1k+2CYq6KyvAX6Q7W1uSDoOxu97SgBvqwbEIAbjiiPVAKc4IV2FYFir
eoSAQg2RGInSONV+yvFaQ01Q7h+SANbgMmSI0c1qCym4q8CF+g1IMS1CSUmdw0CSgUkac9UDUCLZ
bfSUXLEHXV3EI5UyOz1v//ePGLFCZLSxfgkLd4WNm5GeHSn+5LNXhTXW9xDHt+ZVpK2zGUv792ro
A+huJ9ZoUrVeOm8HLBegNNq2coBaIBTmoY73gkZAZHO92CjnCqrknseJ8oz6xSpVvVNRzEO7A1Sq
5daSfMZmPDamfi4ICPrVDHzxsm3gpxnyho47LM7V4jSsn4+i7oEWlWnw6DrVjvQHShjSBN8lpeR0
sLdD1L+R7iBnHuRDAFX2Qbqg75ggigTnLNOeKdb5UrkOQeln+TTcaTM0g9guqmV0XWWHsKUlpfVo
gvZ2DHfjEdEvAUWj6wNv3VxvjbztlK+31btyooBlgSadh+wspqyiLFJa9PieW6sllzxx5CCNTTB5
EHfCPu4lo+7plewapNvxe9rH7COhKOu7TXUPMmlfGbU7FfkRFVgMIeYSgw+FJArNfseC6G27zgKn
UA8T+kUz9zlNLqZQtiW8JhmqnuUiGszLZsLI+g+PWZuff55Dyeo+GmI2uqnnI/Aid0Kq5uS3buBO
VlYL1rVnQwk0Cpr4Xtimr6cH/5qg8bgN7G233pX0g3r3/10U64HZveAM9sVas4cc9S8q1t+Tj2qg
W90ZxnlnyAKsFdPMfnTTWEPTQo/8JMO0tGe3d6s3Uz+Dja1xF7IWsqZjQxAVLuIzmGE4NUSO7KFe
zmNqfGWAh8oMHVCiHd+9OOCJwNqSbKnKOsaKvclS1+OE3Pb6bz/3noPqw71+GxBXtUVep1tw0dT0
FK5JFtcG6zj3Zai+R3qHKreyApiKCZdC2u4gAA3eonZ4Q99Fa1HCSgSqRMBtUjjrOBKuEAfl1Z0+
2uerKg9c4UE0Wi8pEP4pifonbWar23RILFPWV2IMR+hvcndMoOo2S1xzE1k4mLSlW64xbtZJb93c
/E0Itlk6tEvgj1GGyK7eNiN3LNvaH3xiFccPqJI+22Pl7EZI62Pz9RX4v9K+rlv6b37TTa7xQ3GE
bDnkBDrjuAGhmbCiOFUzwYaQUl7F1nIfCLDerw5Go4AAcn2C5RGpzmSogBkgMMe/BEh8htB6VXL2
QcSjH6CSSy3CldzbeD26TgYmAbt+6DSMxDgC0zGxbg0v4xBBtAjJUCCdaSOvlvpOtzD3ti1lMa0c
Y3Kx3LtR2+HWwcfphRGwqrwuMfnGvyZBtRQk6yX54AIGAGdN9lPIwGmMpp9Zwm3hsSZkn2idVcHv
l9e0c1G1dbt4FvddtXZ0VGAg+r8AoCbADzdtzgR1xw/7sjwivUw3noPIPiUKfBM2d5K7B17kMcP0
frGwec36S1TzrG4ri6ttIp2Ahkm0TA/oxIV3lHI900IhDWfd/erNnng/hmrcBYBePxUm8ylh3Nc8
8tEHl0cNDOnj62ce2UFSehICQ1+dKr8wUfKkjRz7VyvQzsZsbiD/rSmCR5/eczQ3dRjpu/aiv5a5
fCSURHAuVZRL3q6N9+dtm2ujmo24RDM3j/emNXJjjLiEsEdQNVvPoT3oRR8XP6yrF89f857+5+yH
oZJZ4pxtpcj/lgALGFrF7AuDxRrQAkcfkn4YiCzYMVoOZYYNcYnvGFK4KT4tpp8lAHnudglz6rKn
5QDQe/OaFOntC34XmJXQKhU3mn3phWZxI64IoBPvWaq9MQ96RjKl1yfTNWDJz3NLIYWCaPed8fAc
mtmx/VtPZ93DLC1lUtxta3m1ImX4GRs3V0OSoJTdaIE3JTagURoPjEPK9LBHuXJlfBLEfnoQ89Ff
Jg3v3WHle0SLUBTymzvUjaAtgtV2Nwvc4anme/E/yVON5ymX9kuOM34K8VlciQDXgehSlGFU5Tuf
o/5oW1bh/VApJpBJBGV7ebxjDKP27wcl6l8iDk6epWjaCxTQBtoxUjlVOrBHbfh5MLz8cMzfqssY
H5IIGGVs2oogIwi9Nq5mxRmGXPgKsOCnKHMFkr5NJq/+bDag+iZsj82A/zCrvpdUWE8jCuvC8/Bj
HwsC5EdWDx04dSTHfSk0d4DOYpo0ugTiiMnH79tT0aiE03RfyPXmTuxXrPTTNrctoBlgslrSrqqh
5IG5gwI1XiQBrDIsTtCqLNCY9WRMntJFpCVPJnqDR2sp4Prz+2i95LlG77jFBpRY2YHMe3JUIb/f
lIIRi8558ogWuq+iLRPeAQDQi9KESO7X2JHjoP3hxjw8Pejut0Ik8ydvb7cWmMaqU09KX3Wclbhl
jWhxkzzj2k72TyAYTGg1Nu4NLIx+VMWHLby385MCp8cPu5W80ixvjQbrfJmKT88YgcYPUGl2z+oA
pZkLZXrcjqCb2OgQ+kj8ak7gEfBf9R7we3N82pk2n3imgxZYiSR74ZDvtmq83uQcMC2ZlH1u6Ajm
lRFnklmQhIVgqhEzy5Ir/ry+HzffgpR/qVFM8Umbd2HOn+p6VThW1riBN/HUMXG46nCX3OU+A0/C
S/2BN9PTv8oaG2m0qwWE/8s56t50KJJYyIZGGerrXMoffQ1xBU3G1MkD0iDW7k//Ak68Rjhy0YxE
yMcVq0CnbMIAi9GqDknLk/wHo6ceMFoNKUHYSB+U53tggT4Ciq+lrhnug/ZvxCrIUyuUtmMRf8PT
Lwjb35ARpgi/lZaM4HdYh8G35l8lWx47DVqwqv7CFclh7WzaWtUeFYwMc9GMM5g1A2BL/IFJ+Tuv
V07d9WQxaGy4RSh5qqKJgT9m7QzpnQcGrHXRWbQ9K0DCSSiiOmrfoCNY7uhpcqAWV7xp5SFeNtfX
FMYHEokYlYWBwxUuusJ8SCLRGmaGuED2bcOnOX0P1vg28jzcftrMQaHVDwdWa6B6KSxDpzIG3zzR
5UEpBlcBRav+ysCOCvbww4MQ1ESH8HIvtBck7TD6m0y7LDDmvnjVekXCawQmNwMuGB5u/a8gF2/a
A9UzAjEHh3tFdxbl3z6ZdoI6xrmRXS4p5zKi3lEz9hT6TjZuEVKYVjfs8iBd+Zr0pisHfpJenF8r
JcKVQHSZabmUaOom4NGzZcKF3ebDo9zNQ8ZVv0+7QUAj8CLHTqkAdhpK3l3eBNGKj4mKpnQKXkUk
8P4/OHa/R1BYB+8fM7Q429Fast0tfIn4l7pcX1UZfQJln/CtajV05IUxj8yfm44iMc5sPv03k8W9
SSPYn7yBpob9Zf3Ds9QIThznmYrOAKq8quj5fOZIdKr9reFSaUkbkumPZkqerlVOsKfRTpZ8mSri
PLIfW9NAnaGeldBNAmNTC7VClooOKJ0nskD8gHG8Qa5LWMfUYaS4xfUVHCvstDa/fjSNfpGsvvFV
8JXpn/+4h/aNJ0jAzmEH7Lr+Hr6s9HzQYghOuY//db+0eYdQbIv4/q5Q2TIu1mnHyiXGbVvWil8Z
UbVIra4zg7muC8pJpmgjNQwr3hyA9NrAeHAQJasZhY4/ZJRx2umLo1CIbDuPj6XFzt5w536LblSD
2arb70Dp68yTCQjA2+HtKZlcif0V1CUhudgcaZQ6IXpEJtNWCeNILk9YmGsf/Tv6pSZokLv3huYB
5vW6WusgFj9Gvpe3wncUUKqHVs1LfdKwqgkr/uaFJ8jf1MDnG4j4F4WyWMV1yj9QBZZrkhaaYBHB
ghWIqTTyjJBdQUAZRDwZutT5faQuDGwBvgDalrrRtTOtu+BhZhydSgBDVNUD7Gf1iieRcm0RRwGb
XhkQoCFiruVuF+4pfMt5vd33b4i+0sNajGUNBJVEHz22b6zWV+Msy11OeljocpgaCkF6O5qC9oSm
Deyz6Em5FfxyGbEzQRvkJoDIaM84iPd+nPqL17lmVDB9kpBN2u/lU9V8AbLDvoR4Dbmm1kvrj8ji
Qd7A6j7ELSpk4JggY0WmMN4fDM1bB1ZO9QatdUBpSaJnAF8Eg+UWC91cFiJLIYEeYkgFuJK1CgBj
9LRn/tcimY4KzBNWA78tzTOgDDRWkqHhfTgOl0D+fGvQH1/YtdNahg6wpyDJrPSzf3omeJ9/wMfq
87Lx4dAgtMNfVBB/zKRWeWL2SjR92J6eQlKFzYFhQL/PH4Gvp6JyC/nd5+SzuxglnWooJnkZAu/b
OuxwYJW3NfgZuUCJz2dHwSSV0dulsRN7oY4TCq8d55DJTG8JIfBra1fFdbDvQKvdT5NRRGYPTCWF
kXxi3TwA7mVz0SOSWTlWgX3JlSZMSLUEJoVQLrUs3BFAeW+rk0FECV81nsiqk2vBFKdQ3pn3OZRk
J+WDzl3lDid2+0uVR5uoTBaHjmXZ7/SHu+g5CE4bVqdDXAPb6KWxxNizF3WWZPiFOVtW0gYXvEEK
trd6pzk3cD3x/tRbdzCD9QACXAmFPzA84rz8YQGga6NSEMuzf9Q4RrOmiC8lunwGmDfYKOGc9pHJ
b0Cv2VsouivDCCwQtYoue2BkyaITkcFzkq60ylH7zD2RfL5W48sZyUESSbRiWFvmBDY/24211iPJ
a8/kj0HktekbeCTVIDFtTbJjaFba4ViHYlgJc4SOrTWyFkxklpsgF5gSPjxK3hFEdoYzIoAWI7e7
Z5dv+GRaKdsN1/BnDIoj6H7thOTjmA9HOeMuzG26TQnOPTYhpe/Ge2U14CvNGnz+tOGIo3whqMd0
IrjbmGt4kaGFRoUTzG+p2XDndw6FDxhKPsxGMj6KN7PX5eQbPeal6QQ880vfM3zQFvkitp6rp3PX
zEj/LDsNXjNFgCa8C3EBAMeOmQMvvCFiV3hmuyXIHWF2nNgIaxMV06oPKcq16yBcxY4jCSR65Upe
uvruTnUa3YYzb0GZNiVs8buKsJMTS7kx8i9+cBodwI4tcn8NV72dHEMSQeMAPWXazhERtmDuYMHC
UbMXXgLTKHVuItMuqVcBPDidC79fYeKWL/Sq2wWMxz3mpz7U0GzBrgsbLE2Izzady+bdZrjcFjmJ
acUo59Fke2lIQThmSM0El/li3W5w9hx7md20rAzX7hEweM383WVaDpjFPvRLeaWEmkdvWXvBbE5G
mBXqGi2TussSwd+LYcr82nKE9p8/ETSaoTosE3KLgFjTSYARo8PLa0h5hF0pggl6AkJfebepPmWA
i4LuJzmoUr5wzgQKfTX96vsaAtv7ImvwwLJog3bw8zUtcTS8AXzh72NapBp9RRbsVZYvqZMBiQkn
2lL52jyfJPvUEoL/Tm/yJzcCDvhJgXjMe9Z7fShLWXeGEKMp/dC0DFKzcqi9Fi8FDwISdffcKhLW
H9xgsNMT8b02fgpRWV92ClioJjQLajdw0Ok8I7XnPBLFAJrc30AYQxyOvS+wN1Dos6fVYhHMZ7L4
aw2kdXxt5g0+EykMpn5Fqtdwg4D7hsa4fJm+MTWR/DFgtBeqTdqDJ/4zHsr5fSiGzb4XYYAmldhR
mjBDPsgMQ7fyaihuluPcc0gYfYaDlpCpp/jaseh49P5GVe8edmPT6movvuw3Co4Ce5qEpy8VBrBS
Oj+IrGaRv8INY01ZKCQmQHtkn+S1k1NfXQq8V11dl6k5W9uYY/91o+ffwwpmhYzR2b1aXkaY+xGY
YUq6V3EBGoENBDaZkVghqYQuvvXyt+EUm8hRE228HVTXZrZY2pEfpm6mn6RV/JlXZIASEthnMtcR
hoJtgzRz8UNJsz8DcSNetxieGiBbQP2p/NnbcrtAJZzMx70WrvGvAGIzfkGUbRhCTqPfsxIshvbV
OGQtf2BUoEiQZFJD4sTOlzQ0ySbMWz7Bs/1ZI8eU1PLgi1l0RoXPCNbmHcXNclxPtVj4o1+wQ7gD
5gePmKQt+F7IZbJwqcJ1VPwyGWlCTMRTZtyEXbzrL+bfTZWiF/qrjLUc3TPeSxCpx/kbqh9hOWq9
rIzQDvdNUqoyNiUA/bFIBAfPjT5PD9p1+VzPDnypw6pLb7eckAIYzI1jBSf0XjRgdP76AUNSPG0o
Roc/m1K/6WBy40aQ964NYRkVPNb2JCfm+CZ7PG+D7nqTQhxnmyamd4n280mRH3VpgZFgzcKFONuw
2jQjhn8JxdUp/wGNdrjq6SAEC3mfncl2960q9ybnYQhpT2KOkh5r2kZDssMism2cXDhlyZASvfL7
KzqGZppSNUzCXIBhfg+l+kzjRZZLiNMXWUT15x9ISNATqgpNYKbqLLDU6F5Xq98bv563L6MdyDpe
IzBRqEh24wkci9hCuSWKD8E+RPJDoxKQ1DTPkT1zUjN3LLlr6RCPZEvTV8/UDwdyHl9zmMhOQaEq
YYMOBeWZLBYrlSfLHOtvOLEQSbaqZVlqa2sz7pHR8UVYhMNwXqEQXkwEvdwRq1feMc53tLSwFBEz
0m4qWmSoR5n2Z64+LyCQz1F54i8WEJUET/NCG62wGplu1vkajr2I01HiaC+wHvlHUkvPFUpV4EAc
Q7Wf1HfoV771dyKDwwXN2nRr6F5kGQ+rx8/V6v04ScgrYiiTm/FrNhzILiftZHtiKGI1Wsxxu6bE
pSzDJXCReYJVRD/NvgddyIYJGuL1VPOfZ2vaKicHS1fdUjmoZQEhPb/D+VQ5nckx5pY4prCVmIfK
zBDYwjk45bqJMYrmfzdFzUlTCDZTCaMTn/cm0Mk6dO/xjGE+10FfOSuZ7LfdO2f2H7IljVzTg9MC
0mRoad3YUzI+n4xhcOT9TQZk1MafW9M6H65hLMMF4j56ZKTE/JCLUAgE8pL7riLB90R4e+QstGlO
vJsevpvfAf+foPQf7+NhqIaX+Nx0fv3KscN8D0YuY6ZPL7F5awGyrjipze51GZEbrbkoliCrmPeO
1PqqtiQpkDUtEssACfynMHpseMoLZNqqasRr3BKxnSG3ArnA13ZbvvQtjvOuWZxzOeMeeM3J+2G5
eRes+o1QPLkia9eEqjH+J4UNBVzBd2SPmI3EmCQW7jGOMPjrvE19Om3gyNSVmvhlvlbZLuFamMTL
ZzMpQajvXzZ3UmtV6vU9yOcNtm9zqS7KGoFxNnXF53wn4lFV+HwG4VsCOzK/L/soMUrv1u7SBWgP
WY4JykE+SkPJdAp3lANdMz/rV0PQJ+NuVSgn3eYRWKBf5hx7qxhSaMx2frZsKEITubEzvCXNquvp
JpoTuzK6GqTb2tIxVAbvnqgh+sLqG+0n4QnKV1RAsf4lDJlD1seObhHOKaoI/FZ6PNd5lF+SlowK
XituF5HYi7LbU2Sl51QV7+iGogmNcpA0Ihqz62JLARgoDXaATsROJXw44tQcp0Ci8n6Ftcq0K5BI
l7lB9gF2jzQ6IK1NnMcMJLQAds2DGcxdXhQ/Bj/4MTucoZ/+DsjR0GfH7Zt6ES8pun464MWFUvuO
OOyI3aPTVfhZBr3aAdRT8SBBq5+d3XvG1mk+qZYHj4czKg7hoAvN3RPeWqD0weLCmd8gVwK1K8Wk
OuxzYC39khqm9Z3D9A5J7hTYjOiFOH4bqQb/bhmAxfWelgCTPJ9CuIA+ww1qCtqdCgZjVhSQV+w+
49MOZxoshJTZXnrWecP8ljD7IedLPxvJ1SzIS7dz0sLTEhAXNbP0i0ePe2C3iyQYq+mzUw3hG4vs
yjxp1uI5MMMLcO0Tkg5wW3cOJLyq9MrbcmcGXvDg96rwgwN7gQABfVhfjGA0saWOoXOXO1nNCubW
EJEpILUctXC5n9+iPlsQx3+5+cIQ8nTM7Rrgg9UmdvbDZD6N5yIWOoFBPokjWp29Urk3MPbIKX/Z
n4pWEoUneDxQaXQTPbxrUUYk+qTxixlZHHoiDeObBrMbeLxw4NQ8oErWHiGN0eyg8TWrm3zsrbOA
97D1Bv9OgYywqPQ4L/EaB+fsoc3uerJ3vAn6eBuHYyjHVM+JpWz3LMu4ZyY0CihrwTrhvMmkZF7c
mrJ7iX97uDGgBAmE9MObhob3rkczjEr5KAFfkMuhsX5sOOBRl38TjJn/70UffZm3O8jc8kGotR2f
aXCA3RIx82YFMSzOFYmaQcZvnL1UgzBfpz9OyycqYx5SV2sqU+jTIyzXX7ZM/QRbGVsJj6baL+DR
5z5j7phcQ4+7uVyF3Y+Xa8CQabuBAWUh/d0yms/XTcz7LovtFrDrRyTm0RjrGdJTrMZtbKwJaK3f
mGvD5HB7WxQwgxDgXEgE1ybZv2WdP8AGhQ9mWEvHbj0zfTY+/bzhAmoG50qoBnC4R70p84fHuRZX
Xz0hWW2Jmj1Puf+tAJIoPMd6rJSGE+nzOdRJfOOXcjuU6MUkdMqw1jR1PNZ04/mGJ0u1cMZBszpN
UV1bqeHDxoQi3yoBotXeHQ0Gt2zrN+jJ2ralVasAeJWRZUydMSPA1Y8Oc+1WZQgPdrahLsZQUHKh
FZgYlt0tDfHaxKjDhUR6l2Rm+cNhdQQmEr5MhOhTkgkBCJTdYMlkEG5jG6vzpEp673W85YwXfExK
xN8ZmbMVV/HCW3xsXs0T3bpgYf8PZGURaDbOc1kMVBp0XLmuSoFx/jstbSeaWj5GHPxJqnfdpwoW
M44QLfdbT4A46Uw+nYmRyi8Hb9phT7dajFXSW1e8XAkvkvZwH2TCDF+16taiVliOBTbViLZbnoFj
rw7MfHBAAVHj3HeVbWM40ET/QOL+uVz3zl/ABTPg4yzkACY4BsqkK3yjarQN+KljrPVun8r3FZAm
xYuLlfJTg6oH9P9l/+sgTsUQ6PxMOcnCIBdyqBgm33PBW+MA2xqVtOJKw+lb1V13eRFACY10fVsD
VwUnz3WupiIT37y01FfIw2bu8TN7lrQlCkBdPKvw6hXwrdUVLB5FDc6RidA79O/2fyxk8hvBEt4W
IbHzPsd2kQ/kDxBWfZDAz6fZ5Xf44d3B9LuOyRYdNR0Sn6JPov4lW6bZC9ZGvWpKOOxdbNznIj/x
RnxV/40lUOJ6W4PB2AG4Y/+Ps0ZvgTfjAE8zaz4LLLo8ohpO6s2N5ktrqcqYhb/K2dIcr0MfLT9a
EgfaKlzxXKZmSBdSjU7IIAR08ZWeCNCqbn0Rq4hJ2Yt1zz3WfSk9aMYDMHF9/rxBHwaIluWqw6xF
vgsA9/F4mfIjefrF+/ZB1DVvuWIG++5xccH+4e3xFZNb7KkH9Lr2n2w1EZW5g+0IftINdltuygRr
04hGrwat6Y8aNHphXvaAx9qZuse5qhpLUlei8PnkX46r7jzWBPq0hi5dbUWJhHDQF+cI2vMjJGc4
bF6PBTtVDNCcSEMLGJ9FaqG8/9Xg2jRSTY2C16xROWlUf5npHXLK6oloaBO2IcNJdWS7DGC8KsCc
LD318RO7bRe8w0TjAwrRYcs6C6B2abGZFHxKTnjaFVeiUro5ziTcNe/jAKBXFVzMtsHjC0w33HIN
gmtYYRiQP364jJlRq4uq9grxV2X+Nct4LapdwEO+xaQaAtJq/ck86u/K46nH0drwlSJTxINXMaVJ
kMH26Eg4P0h5MVBJY20qFQghy4XjIBz9r2aiRMPjK39Fbl2JKHu1dCQ8MvSszjX7mySQAsvj7K7y
L3uH9/a5lr9K9o8j80sccjvRyo8c2oXdl6//8b3aAVwPtOGOpxFIxAxw/B1ot04r7afvPcV4f6EE
6jOH6iPOUrB+ItFxuOQUfbee++QvdN6q9x7xzcbLo+Di3kZR7ywGzllRZsWsdMLiDl3s+T1B+ytH
OoWqgPSZ62qJ2H17orD6a5+Jvu3n+BQpFvjDxkLGTIyovEGBh5oJ6IGS+TLnruPiD5hvOQeo0TLb
851fd6sP9lZEq22H0BDHyE0imAdx4SodnGLu9MCRozmcVsZt91aLXWkiUrtZHEyN3nmnSdEv4ZsA
Bc2hkFBa8tVCRlqYW4xw1VUQzT4FK84wAgE50BBsFLCMCT4LX6LnqmhhdEjDL6e7ZJn6CwxRZNEY
wpUx3cW7aE+G4NtZXf5mvo8RsULGMGkEyUpdp7JFjqntU08wzzMEO/jjbsNUuGcM6uTGjt2qAyUG
356FzS0p2gAPmqU8VX6KShHIkfVA1rYhHrFG2n8atLN+PGnIBQz04eh3syF4NUlJB0ddS7Zp0wx9
R9EPZZ+1mF+FXzvsvL611uOFma7aT6rz1v0nZVsZaPUIBfc+J1hd+s8hOZ/I2WKx78p9yrQiSUXr
Pna8wm/W9dPAu8yKW7VpeXpMZ3t5D3J8O3QArfop1ZaS4iNnvIqEaQO3AKmcG+7HImkuiJQvQ8RN
Brq2cYleWF7lm50PpRCbMoCIEcuED6B/h+Ph+PIKRo+q+K3UkfMcb/tB9Dn6kllSzfOmfuGuH03U
ykzs2P/oZhhdwaWbox5H67tsg8GNj22PLtfT6gIIztS3QyVsHkjihAZJcSeSX0sHo9mSnqMzY5e2
djNVFp/Gt1eKZNxmvle/cmWH8Y193WMX7EOfUDOrMu3PoIGOvcvkxn4IcSWHm7kJr/gdKmhrOyxb
ituF6OcTbK+AYClsaPnvUYikt7Ych3XZ3nTxrugQd16bTdkFrN3FT6GMrCDAM4C2CtYx+U8jkMWK
qYulrpWE+LwVnNAEtOBEmgwqcoecliHurewdz5qdi052unsB3fekSd1A7k/fJUD5y/adTcsjMPPS
E5Fv22c5WY3c2n4o/5HmNFaUJpGlNbXgpaq6W1cAO9dDJDTbGGFp9FgYgfbQTvwKiwC1/ZIy/6PT
N8T44Xd/uf1WA5ul7f4Fl/g8zfH7ch0eVVYX94dU8vP+CQOzM/WRYOfpIbEtO1Vvrj/h1gonLoFo
JEE22sv3gyZsAwMcvxx/K81mexNDAn4TGEHS95D7Asz3U1deACzcf3stEI6HMEv5Smg0EQWY7MHT
mhwh9TemeFEdr79S++Fgb7N1Pwb3juDgz5lVKo32UMjR6A0mCiTmD6q0w7JYyh44KA+mxKY/7Ij4
gapSNc/EG+m0UiWMzt7tp7eV1cVYfuCa35CMQtkGd5anM8EpHhSoZx7KNPrnd3C6kM8YZO+aZFcN
GFbigDNvbJdT8vpQ9l6gtER/NVeBqgJgx2BRFa8FAa6Z2juaGyDtVjljrD8Tjuy604QjNbyeYEYj
Wr4+K9UidVcHUqjAutLIgvs1ltQcZyeLc2VwY4zLZD6/4665/0Jy4VJUnQ1Dv5XEbUBhSL8vEwel
tBSBnKaVfi3bbMcOyVFGQtRVhc9dC7ZY+Me5rdqcEbzzCX2TNCb74Tsvo/gTf1dBg9lW5hpeti1b
Dsbqvi010IzhaC/0vAp4M3nxT2z3Y9UxT9O5sLa+udClQzIs5PZnGW5Pgrl0lKn3N6lb4luLje8L
sfMKNP7cgKb0PaZjXidn+gdwAKeOGu2UPirE2ftSg5ziJCTOIFueX4I+7sdIcXJuo50wFlM8YWEb
mOLAJGiGK/brEpcMP4EOenRjP9eGAOXZcsZMZ4sP8lNNisjy4PAOyb9edc9gtCYWJbgKQTVgx7XQ
Dv2C2Gj3ajT9zk4iEWzV4AlHt1rCS5qhXQxbaGAYz9BtwEVFnwpydxKl8cP8gmUTITxey/iexRYd
WQpETklTxNpPFxUxcKjTS+BwrSX1spGf54SVz57QXbFxM0f3ENpOSyiXR2s9rhgcaliYlO+pFY7I
y8J3Ek/mbg9jAeX0JHB+VAb0LQVuRSwwbezowkPyYgdvyYI0i3GSPO+7eVEni1fyQHUpVt+3L5HG
bg//E8/fAW2mLkNQPmL1aaPawCExECjQFW4BthgZ6Xn/JvOXs1EHOXg7WMvDsX9Lw8jXZ8wfPtQm
bwbt7cE3neQNLHMNxjUvWhKiKGtfQv3Ci8bw0BuTusItmgUID/FfHG48n6kzRkwW9OenDcNoT9/V
ta85mDEvXGX5Qr2YQJhu3m7wJJODGdzKqG2Se5xuZ5RBkFiOwCKRHANXdXMdutm1rlLYbpaGHY3u
tl+8MXsBt1Ud4SOqXNSgusYK2Op7u6xKfko7IoORhURlpMkOm2jmNxZ37jir7631NFgTpn/7PHLT
accGDH2GkXuH3POGzuwLNDIgBBH35w+89KYtahG9n/3YBgMNnPy/s4ibo6kc3rPPHVyAgdGFmJfc
znOUo6W75dOczBSd5BECh0oUFrWDJC79iICfHA7xSJ8an7zI3xNmB4UJKPpsgySHrJlYc0UVODUw
h2XGy0U31PA1wp74Ly2m3akMObeoGCYx3RNR3zciDTZdDGjwQpvsmhRT0lVPL1MDLRCx1/UCJt4U
kiEoTBIxWrjFApAwkjy1k1D/lhzewDGcfXDohjzNB0tyB5TekacUaUUX8UpRADCdeawHB/5VcchE
X2Sk3hSPT1C9aA3i8LVfF8TuekA3Tn7KcO25K/op9YZe62FjJflsZyZbHfA2LAL91GOdFAiC1NTv
Xu4YHmF0RhGQ9nHN1RtjtMGimMluceBQecN3DiSJEomkVeJ2szSMqaKx+cPC3jWvJ/MkaCpyYAzO
apuHBVILW99luM+7VvE7+Yx+ZH/+PalETFcYOl/Sw5HW+U8daSptkefzbhTxtam42OK/cOxylaiq
LHUAahsF2R8kuT8/ggBzaezUKPbjBmkNPqAyFiSrviciFMWW2e2CYIIQ/kg1ra9/d+TZexaBLvyt
AvKgDqZse1iJ0k8jiUvt8NTaPJeFuL3YA6kQ+QuAVtTAI0Bcxpji8sadpeETMQOwkfVyjsRKIDIz
zX8ttZliUi9jvgFT0XemxmTIve5WtwXRtOAW7z4bC2sOn9mMHoy9zGSmfL4cSC8xbcsCxppYzaxd
YUXhWF/HBEfl16tQ1fmkCx/FJW28e5zcQ3ukr8yjwZociimR9E3BMcxa1MzzXiYbI1M7CSgFhJCa
4M+hKuDHiNwXVFcUyP+A8Pv2k4iVH0lR4C4NDvxlSsCzKjmioURg33OS3lyedxa+y1x5zn5pBKK0
pJccW6cGXrd34hrUgL3+rmQ22MDAR+tjkeh12Oe+czf89IMMJrkInmwkpUcsFqVmCHonjqjm4UrR
GWq5p564/l4eHAu5aD69LGYqIMy88TiX/4nCXxk7j9y2rHqHORzep8GhoGavYqGqZ1fpNDIJWqrt
gXkgJpFPW87yemwon1YDGmXOsH3ATPkjVK8DNdAwO05zOJ/dKru7dLowHRHlOOmhqoGKOJ8a5Rjj
LAyX1mqYL5HT21nwIXUgMP/X4fVyjaExFofRhY13NETmfKbp6rSpxuPPWPssAEjGkevgHe7T9ZAm
XjYjL//H1OQGUF0fp7xba4vntJPuROoaBxu+1PyoRXIK0Qdrw8kgCBjL54YR23uHjadcEuNSiKMc
0Amkh93mCcuUG0V/yzzSSXk7bQzxEJ195TzvReIyHf+6zbs2MTcbtvMbS3Jed7m4sxOp1NFMXH9N
ZtwiZEPfppuWHsc1RcYYRuTYbTZNbMDudVXutmtffiaKS5f5exHN+gJf/v/4c2vPO2tcipaNYaKG
SBnkrmw8Iqx3RU4fbiIxY1zvgYX4Nz5sDl4lOvp1VhkJHX4GTZOD3TpvMVwUphGwRLFqgOwKjSWv
i+5ER3LtpyH3K+61wCafHUr1R1xgbYeLa1kwvt0eWAK1HRhFc4RlSK4t/Ccw1Dk3EvtF1uaS5Sw/
DGm9MwYSP1s+g2KKlN1zopbN8JYv8fq+YDYTXX+xNG4YX58z6OsQhmhN+xGm9EuK5coL3KtFktns
UsaMzrmVhA/rzFnD5JYN91+OadyOwqvQNS/+at5qFENf/xxSGWb9QoD8cxsiHnC2PQI5Bl06g8gS
WFUyD/2hItg1FYkNMeCEU31uFfVXUK7EcBpH1FhdPrudr4v+3B7BhdNB4pHAXJzNYrg16EuqD8/I
+MCTeni86bejw71Stw0QHXnuASwgh8Zfly4Tkc2rJeRwq6tqCcJaJRlvudpkEN9WqumcLHlA1Uls
2Galk35I05RWDbdDogjLczXuXubgo2KgwbqjG/bdcFkHVyVDO4fOMm6k87RdWOzZfG+rx4TnJ7T7
MrfwBgjIAOdfKc9eKTk7tDA/KC9j9AX53e7yiXELSkeIlBZUj0zhDBLwJV95k4qwmV/ATwHLPJ83
5/cH8cO4u7UwZJlkFbqVth+BPFwYQ+n2rNO6g53FHn7F8vI7I4HuWxG5aidj8miu6wLa6rcaD/KA
I0e7KTAt3IRuZyDMVTP27nFhZ3u3Ez4u7sByHQjpsTIhtqE+neh5z98WzEeakV9jBBNOvuEm1n6T
KlzzZGeFm5sKm1yvvNKc3biNuMshJZ75RLN5cZ/kGEoiIyZZJTWS2nsRk0uLfAxUXt6krW3fkQye
j6iOUZQbk4KyTSr2WygZ3xBXqhXUSe15I786tGMUKpzUgylussHqv8voDCp9mRp/ICbWkrDHbf7l
FuG9fFsmZjEfS9UOpuQYtV0jwzQWkVjhzkBcIB6HnozWJGg+J8OCSC4H52HPF+6KR0jgHfH8fu6C
Cyb9U3W53gKs6nh556OpLJZ7tdiPmXvX5wEF9A004XBDSasypiuPqBcc8NG9PHB7ckBihXYLWgZd
pX5LD6/m9ESH1C6ye7xXjHQEO4/yAT5ed++efwQPzi/QIeLAZejzFfyE2LgQBGqa+ngT2u5fWXyI
QtTxRXiuWPr1msaTKkM1bFbgqiKbOj0dTyqIPaAcY7WOoufxTrMlrtKSaAaPhuqu0ZXPmOMXS+aO
/zJm5x/7/e9v5HuqnmwerCIMX2HwU8u4pfrTtNHQBbEHrqSkIRd4GD06/qwY2D2xzqQ1AuvKCIc3
tdV1lwzPSxSgI25s5T7BUa80+fnD28BzBjz91nkTI1J+1b6d+D1jdgUV8ntMjAJwE817lgkQKXMK
/K4bWcPmREe2eIOXJKLnR1aAbK/UBPplFWQgqw1HvCGVcCVxaBBTC3QIcMt/cztEyovVY23jsqJC
I1n7cWOsXYkUrEXI+knJ09Kw2JhO7fV1mW7S64/88CdTuEmWrF5hnLgmCp5lEdnxZqnFd4QoCRNZ
ESR1k922xZKl8QLsg87XL3nl7Yhgisa9EXYCUHCRlyJWtZyYViNTBwQxDFMl6Y2wAfPYysVSC9cT
Xu+ta5Q5e41UzaOZjOKh11vrBWVC7GM3dd0mbPG306CHyhfK9gmzRdXhMSdZckZESjnibZaBbXAH
cQ6EodfzBTGt0vifNgZSaN5k+++KWdf6iREzy67Errekw6q69l6jmX8X7ykUaoutaOIMfkckdsBx
x8IJfwSB8M8xTH6ol+7QcZ5fX5J/q8NXC+dI69a+1fXxxYEjOEuBH2PFHccT9jhBsLUKBfhOvMAh
qEj0MBJyjyvfoxCLPLySeGdXMqyOxhDgiI7WWvjXzGMgfEFPdykw0/H8kuTQVW5xIyzmk0cXiSiw
+z+5mgYC41kPyaf4X0lrIuRggfPjm/HC8Zp/Ez5BY05KiI8b1vHlcb+XHNf5m2VXhDwz2+ie1+qH
OqnojjqhhmbsbETYLOInp5UV+0lEC2ZybHUZFS7kx0O/pHeKKlhXoOppt6uEZ7YHcbuE5yUvgN9h
lWIEGh8OuSKHQFZuWWsf660BTkPMBdk8NMAXqw/Fng/gvLkypA0ZfHnGo5tPZ74nblCN4PuY3HBe
A6CkNf4wGzxTaVxa3M9dw0+2GuR+IIGNyrqDjiGYyfcMixG0k6YNkEBjG/RU9O6EaS05g+jPYRft
RaiVYYErYr0rjBWPodjfaV/c9r6Ezp8rmG8VL92B8UEfQZx06nWNl588HSOP4T4nXxbqT6/Crmnn
+6HBNSOeDnZMoJjRGHb2AO+I+kmapPUQF5hMjHKV1gNqxonFpy2TdIlGyhIU8tE8SmyhlxodzbtF
008aFvYq/q6d29jnWwyLCTYKumhi/a0VUun/s+CsbmzYTbSxK7rBZ9/2yqNb/ykwsv3bZFAj1RqU
8JLOgPDJtnlI0lS1091Vw4fcpaAIoL3pOzGuunoH+ASfNb330CEVS9N3GnvasgOh2Vyqq+gAejn2
jhnKU2cxghGROrc1bnbZ+MJpY87Q4zBRKNE+11hmLiugAf1gGJ31+B5TpuHoKVuNom/Rb8KpOgpu
M1HQDBwx7uETsUMLUwnPbkCcC+zDzrABhggqCOuZfEaInD3NMMeYilLnOPireaR3A/XOLfLqFkVA
KqaK6QNR5wSdVUuryjvG43cEjHfWRoS1O4TfBY5gZHhAtacIAsZqronF5TjvsT1h5RpIPn5H/r5r
ZMac5qcaF1FbTrl/6cOUv6gErOb1JG4b8i2neEGlwY+NoC4w2hNh7AOtT6in09eIndB0DW9YrBze
MkKQb2eM8kYkFJ4sDhwlZNki1SDONpldQw6LKVh4cshYM0aZPeSL802Y1qYfoSjKFGxxI5447j3N
5/yM6emU9TWGqCdoBARYIcwQxJ+17SNkJmGhtSZX7YRAAFFffbcVBgLHxTtj4Xfa+dVYdT1IOyQN
RD0pvUpquICp8EqwF+cBcgswjbN6JQiB9O4n5Lfm8VVdv6atJq0rJn/QYsSIfhabfxpk0Xgs9Tbw
YlOiC+1bd8s3DBM5zpkhc8YMSm7qxFgisedEue+NKpmIpfoikmb7WBasVDUrhftoFLu+2k8ID0gr
1TLHiinFNQ+Fk4NQ0EwB8bMyGONRZw86woEx1Pmr8znX5yBntZ1SkO+zuXpj9FkTmea8UaHzE+vF
NPQm4e5ddB1BotZXVeKlV7anEPULc+0zmF7uxp6Pbvah6FbeZ9VL1axn/vlWkmfAEI2OkvgVe1JN
bWWNzfwXkdEYZnZ0pqD313k5l7gi9FxJqUuFb6bK0x7ECtcz6gHUNhq1WyW42rTO835t6Ln28iOA
5n6mkXHC7qX3LjQndDAwxxP9sjbK/ALC+cK5O1OTyOiFMM0b6YblcJq4BaeS+J70ku8/azsmbgKW
ciRVAHESLvIgOh8erMJ1fp1zb7tMS3FBKU1eAy2wRqqZNE1nz/FR20YXVsRPFRAOEHMyq9MiVsJx
tKyL4sdBj3jV3ySEaCRVcnnifE4s4VoS6Wh6O9tnZU6BFpJfcc2E3tyRZ5oQ6qJKM/bHABeXv5/Y
R03Opbc9HZHG/1uUOVDgebOijXZRMYDHGMIkWI2WrmnASwgVdyZNH/URUU7XhxHuwTRaW092U/jA
yZYOdr8Q4/mAnanN9Ty3g1JMAFk+g0HgDzU+ADtVNzx4oW4Qytg7tZiVyaxitFz6Ar7XKFAeeFL6
M/MxJB7V1azaFkf+ZEoDXdZXeGQ0bU6jLDfVKVFPXPV8cynVN5eneVCBds12+/ikDQj68ASeSxWV
NwXR+afR20he3zAVWBUPNFqA6DUBIsK2ncC/GaQeeoLTthRt62rNTQ5GdRbVKxYwPYl8AJxAjo+G
F3LDo8lgoDhhJ8gwJ9Gvqc1w2KcR3p3uxZJ+xRtfvE0K2jd7vyecXcvXf07lchexTxtkdA2RNtA/
M67s+5T6oNTiwNNXSNe9nYNh12xhCftuZj1VAuHAE61CPuBMEf+pQTAEAts2/rBJMsQEI267JLuB
8Lr8JaYFv6p5wZcbO5H/Gi9qIkOIRxbzVmjGB/6p9M2LNrGWW8kWwwkmcsSrCYnKztEIL1U7nA2h
61XuAcQFFIUPG/NDpcETDDZf6uj6jCgGiCsr3HlIpO9QX1Mk+daBwQlaWAupo2HDQIyyPTWuCUbY
MUUNPNmNvIJopGowPbRDZ12WYTM0BaDRowoq1zUuKiPSZccdexeNtvu8Os5m+2PS51kJJSDP9mrI
/PnTlThqitqzehCne6KdswEXTkb3eET0ezWP1hzi3zYp6qpzRH+DEpH0L7gDKSKwmvBPPjraDuoj
ep2eVym3Yb4u8aK6EmkuKvwqjdkJQgg31LuG87CeTqgH6lPYyjzl0xnELTQKYXMIBOSAWH/A/NWZ
FIktJbeG4cYRi5UnvZubmrafGrhq/0VSfPTFlwtEtQUehrld1bnq2KCmQtrOudwWGoaP4S0rqFuR
kd/sPoTipMKIsg4jkLj0F0agIwqsDMbTmE/P+s85Hr31RfpS95EYZOySODrMJQm1J20C/drBYO/9
WeE2rT9T+EjParUtdrwssw/LLLC8mP60zRd+jVovG2sNMaFqWbBgOwNzI6GPUos8nFku4GTj2JgO
XLsW47GN1TFeKBqaU538mKcjknjDEVgkQo/cN/ZbW89IxsNtYTfrVOMST63qFYtj5WcUxqmgHOkB
M2GpCHqq63MDBx5bWBLF0F5Qon/9TH1u2yrjLkd/gEBaI6uLkEgEy4fMt0x5PkwLQ0I6OxJvrdTB
kcpBlyX4uhgFkIf7v7Kcem4qxYlvsbvxnpFIxgj9MD4WFHd3IrTP1xKG+Jc6pN8Owrwpsr4gCf+g
lmou38+0MiGfpkIlhIWq5u9XwotiqZX642G8K/uoCYNqKsQER0o3thnwRjI1NpDRz9F7FFV6DQXN
9j0/FO6XTCTj55TsGWE/uhzOro97Jay4PLJxBgBFkzyMulY7coHm/KkmMyZ3xn4Zq7wl2wrPU6zo
ztonPoLHdhpjaxJguAGFqTuArQSj6b6HHACRA7dpHfMQX3yqEQeFsKEinVorzJXP1Sc2U2/XS6IN
htrMuhcCqowQOjFdYKISFTIQQ+wmQzMbzYWCilXeK6lTyd1plVLaLu0WgjpddrWGRQjpYjFIaCQR
PUCpZa44LaGHsLWbmUMjRMUFKzdqPU39lGsje2s54sLWeL+ieJIM/gszGpfcvwyrapDFB9FzontR
/MoO50hFZo3QQryiF0uDI8y0WdsJzjCiZMU2P2CHoVr8g1uMMRAjWeX/deYAWOpN+Y6Qu2TYlH/K
yeWgJIBfZamWme57P+G22GlCYoRUVRofg00hJPVkUz+VnGl6ntWJnyoGb7vux+FhRxw6SOFBf4kh
TJzyxXARw47IeSLa5w7WCKAqfIB6byf8sWg7g4ntKuEq2Pgg//DhTz8rM349eZGqDeN+OiL7zse+
uHgvTVe1ZB7NiWKSoiWOohE8wXEaRMj0NUDAxHpMFRDsY/T7I9PVlszo6Q0I+VgauWjzmV7oHBcR
Ox3o4Fx3EB42MaUMyiApmUTPITL7pM/+xUANn5e4tttfihb419B72TxMtWy2vBjPYNeN0V5qKgvP
G6GYrJg0pwUQb9cE1t2rZ9sq9a3OC6Ng3Xpn6M6OUSYHBwqu44w4ht9EYsb9pwYLfcxdz/JZN84M
QWSJE/a9UwkWv6uAbaFzZ+FnA+FM8WsouMdColdfOOcSDySuEcucj/+zQtkS0G3KcMhILZESt9Pg
GUJNUQMqtg4ntp6oOdxJuOfwSWVzyfIC0L4Ta6O+3C4xzYViN1XYpe23bFj3THoaLgQSR1GJq/7A
hu1TJfey12XDREqpvHjtfBFg1+aH9/bMai+C1zZ+mcmieooCHDwUjF8TN/psLI3xQrk32TtJQxlK
f93MhMuHeLCe6rrFobwjB43baJ7bxtHi2jxQRVetMmRSLElGBrBtmD/69Fzj0gFur9QbAGJEmN3U
ggjBdvj3zU9r3MNHU+FbYUaVWic2HjlEPv6mMEA06nwzLRos+irGsV5iRzMmXAC3GPUgsjd8YJmW
aN7Nkh/0SC3jx5+C1A+zhHFA93hE8wrp3h99ceog9jYuBALYeGLPSq+xEGpPlxdPHINK77gaOozs
lWQQmUPzTQgwA4swnHJQ90ZptwNsc0CMGBT05lz0VBA1/ioGRgRh+3lMcV9Z7kCOL2e92lhnhhq0
zEtxMzB9E6/3FWsbcK3qtxe/P8VBUxZebSiiAbocPiTGL0xX80ryIHaV93q56PH7TDXERZuEmZbq
9M+BssM7WvCDa3rS5sutY9IB36gfQoZfp+ef48Fj0A+iJgpi8JR79LE+weAoM+nd/10APrab8fRZ
qmXhTKKtn/lMNjYhXrq5dmlZ8BymQWc2QrHh5CjILumV91QrHJuzrrkuqluOctjHX9NSRy88gboL
HGrHJ0DEMDRC1VbdZSb5/s0Jv/m1Y8firf1juEDONmx/rZlqrcHvMRZ7hVlKRbFVRB657T/z17Xz
1B/TjXxo8fjpW+1tC3STth8gILBhUzipXmaCkR6iMhm8+L1VhlmTNK62bpxXe5I7FCl9wCIYpv7P
XK9bbR2jt/2n2s/G0BLcvLUlqJqKpViJPcVkefswJVqOOgYsBuFSUU8Q+wshaXB+10flzMMQF/mv
JE46DQbu+10CljNv1Ib2LNkKu3lsWGwBCz7IMpgc3rCRJwXX4TO9S6KFWYqoAv57BjfV0+2u4Q8s
K60tVQ3je9SJRTsPfg9NROLsaMii4SUnKj2sBKF97FWRiZcOEmK/jtjnhGAyo5u3EPoBlkb81Q+V
88KPdaTpYKy9h63TS9d+dIxHnDLqopFBFt3KEvLFMBkv/L/cFo5d8YN59VR9fiAKiCX1+wij7mx0
yJoJAQixqtYd5Eelym9UdUYFoPmJGvLXubndR+J5e3pOxvdfX5OQSf+adm/8vBRAx6XWhOcsH9YJ
BcgnCJ3AsZy4LbvhIMayFEP/LiLxeM6bRaevE8FST+wm6aw9DHtTHI1QkfV/t4gYxtZCpnVyYFXo
Pmu3hR2XoliYV8CB1rvV3Js4+bE35YGQrIGHa1+HHy6oEJeyDWCVK5JpoPAFAte6Moy3yYOkzzyc
5/Hkax9DZrlHbeM5oPE7bTd9ULbIViC+a45AH0J0HP37zudeVXMtjddkM0zX5M4NFomJsDeXOFQO
5pxSQUf2d36YisoaOtklizzoybVXw1i4fnB9dqCiF3JraHALhf/3vGLQOakrT16pg5egPfiNrGFn
mQgeV8DwkBZe2fYFoPeB5vP3FYhS8KQq4LM/UEn5FIn/LJm//SnYdUFneQxfY+rzUsc6GNiV1y76
03YkCIH0DxnCxATWVC4YgCzssj3ZkYBPrTp71RokB2NOhsyEjW9YOT8AduSQaULuvvGOpZcxDcKH
Oq7w/xFA5yC916bYtRQ6WvuLaQOj9TQfeV9sWwMg2yXcRsP0Jw0sbHYhDUU41SCbBMZ3celeP71q
7sojxJu2WA2pJ79meWkcLEYbDoFEcRD+yYCb9xtNm9TWfdJT4bvowOROwS6SlbfQB0DM2h2SqlNT
vv4sbZpcvn0Vz/tYK08hLLY1netYeLW37VM8jF8iH9tkiR5nPNC+NrsOKqRweUXXPYPrUelDEDrR
Mj8Yq/04Mju2XIUswV5o4P2+TNdHfi2EgndauQa7wXH5mW338zzVYcS3jU71DGNDD8Op0h1pwWdj
86CkR6OL60aUfLYrIgNwHQotYAMNTg+OjAjVu8UzM016kcGMqMwIIjpY/7tpnY8qbXG0vwvxBtZG
5WYD1OCuAyrW6vB90ssjqxHZixDFBZ10Ei2skq8Cz8HeozUwfjNzAIKh+POUqR6WvTfyzuZF3GIV
fGJXbGQ7dqK+7t6V9FYfmozyxD8reNEGyTobLBNAiwzT0akHRmTgRnBuMc1SoF/+H3JuukvDr/5S
ZIzN82hxUqF6cXU/0ay9SZOuJlthzQExZXsjqPsSJl2XlX8YqgPG395pldzFSyYAYx3qmVanfc16
PTqL162rqsHQlJonvQBnmN2pdZGWfjflWE1f3nRpm6XC6t5mJ7Q9dFeS7rJ+31L6Q9dt/dYYhM9/
rP+/W3VVolUpIQm3xrxgDTbB7N6oaBkB7YiyglxYWBQGcAwDCUu8pjrvXHg2b8OG7BhxTAksaPAT
zw5iXdxOGzblZGl1938uOaoL/dTBxQYYfF2OTSwaCR7/8xpdzE695u/PoWS9623bEXa455vioIU1
k8AD1e9MAtXEbM64HwxyIu7FhXo5voOEsExaC2pzn7QowDRxwrHEZcna2P+vmHmilxlHgJG5XLZw
gnnWdItnF382JDqEDex1lBNuDVuWUJbBqsGxeMTSHp3leF426Is6YPjK9w8ovh9240R8qAxpbsjw
zanSKyO+zkaTs15bI+e2lYLY5qyC0qqc4R5pND/LtzA07f8q6tbXIxawiHbxTn5sTres2T75rACZ
02rZ2efrgdKh+LtqwU/f6HyDVM5LHFQbYkP9Nz54z8PPUmXNCyXjiglcYdM8zJeymZwuvLIsv/qq
PLzZvXQnRbDrJBRB06VmLrrjsyKq2d4ZcMwm7qK5v2fXaoxGZ1EjSMt1hR1aCQinUW1ivXK8hULR
pArjqyNZc53uNphTp22z41czMThwsxYHb+/34afNZO4T9PHxCgCTaiZjSzSbYtid9EKPsS8/JQvJ
ML+22KcWGs2dfEldZDKBnu1UbrC4gHkLTZPK8L1oUTrzQv7q6olOKJhQviRloJuqq4My8Qmstu2m
R9/sZklfLeh/8aRczy2zz5hANtrabgudfIDm61kbaXwVmwtBCGe9jQp9yc7E3DEhyT1ftt/9Kmov
RvoWWQWKqLDahlY6NxTmKerw9zetPi77FNDLfPQny4im08H8QmvJHUMbB1vkePDJOIwSU+h5+NDl
y1s+AvawagH7TcHlfLGdZnFLQHD5r+JzVl3ozvzJvw2zAYWStLWBk8e7vXWi+DZnIO5AVq8KdOvI
GGfjTTNeF6c03vkfRFnAQBKzXXfIjOiK3ElmOAkCc7qk465cc7uiQg0m4kdI/yIebjuZSpwyxOCD
LhyzK7mppwRXAzBBcIxvmxFt/fi80zVzcKbiNDJmZBKNL1PE+nGfbnR9m4agB/jk4TcYH9cxapRW
HlaxhxxrU16limqDz2VLnav2aABYbkJ+n45lAVls5Ya0if9j4IM3tteh2H6ptrn3GzRmIWycxygZ
gv6BuqivbqIy+UyMi0HNvd1ny1pfkji069LZBCZyIFgktjqJwVmf/tXMTU/PWv8ynT4bd7xbGL11
lI6z7/Zsf701unG/bZJXBFbwHnCWld0IpPvlELsuanUIMUP16Z7z0x/NMSdb88dlnz2phJ/C9REZ
ETGzCBppooMdJvR2dIvQ3+TweGbzUrS4TFWW0+zf2i4AjluRtU1cOyGi3kCEnsyVFint1nG6pNyK
ZTmQWEQqKtpKP50C7Guvr9PmlNO21kIxoJ13OBfGYlK1WQ3ZDBMeU4d51IdrNQ8VJVJv8w4kQcxh
fUh4qN/ZC2+zJGSKK06nx/8ZCg46i06cjDE4v+1zQIRm/QTXuod+P5F8bUKOe/CiXgy8vmGGb/0H
JA5wVYZLpNbQKpC8YWh2qI6/1GMRFOHr9UN6CgJrhlX3K1AgcFfo0VfX/LS4PS/BR+Siw54eloKk
2D972z9P0lN1iDCgaArQTIN8HNppLzcMgOI8eageFyO0XlBB1lpBEdW9GTtzpajGU0wgmsoieQ0k
3sWntCaGTK1KhnTCzOZ93HYa2gJqwbFlxp/hm4qwgcasSmgszgUuS1hypiXeNsLv3QHa7x8F8OAs
X+LuCHVefMFl237FQJQXR/KTDm37ymGOpAnjdnjFbD8sWuJ6Kj5xczZUnZVGR8it5VwUOy3dKxoV
5No6LXrcZqEBW27LBhFmV8d0sK9aAeTQleOjeOBxNhyjEbLPBpeaQJLSRXF+2ccEHR6phkdxk8vB
lfhNeMyL4w+LAinAISRXXzSGcED8tIdBarceZ/XkhhWokvIf7a4YWUf9cCbpZ+BIg+MPN0XQmYRh
QR8GT0lk5r51pQ3BVe2e6C1safAGokFTYZ0aWN8V2A8rj5EomoiTTVUbpX2xr7WSbwqIUsmr9oG3
7a8buN/sXjAKBecr1MTPuTPVNxw/W4MR5bvG4+ok4bAKyTVp31Ku6ib/Zncgo1oc9bsy8hZ0uuJH
5AGZVC/CZAJ3mndeeaG24ZsEghzvKsc3aJ7uZmY2ZYgGnaWo0b5KLdvI+8mPGJXe1EXnktXisk9b
AL5ZOcqECRDoDYXrUsBYqiFQGIzB5GY6meuZzWLlmPwgdBAGB8zFe6Lai7Mtt6z6Mbt2Y90FsKc2
1H28UMl3dH8jiXGA+4aPqAn/fu0sf+5tzalE1YudKK3F6ZXUsRuMrJqRVbO7wHm5Dr5xFH5mMUYH
jCOelxLDOHp3CcoOPMTnM8AYwVDXNmgUH3FU70MpNeDd3mVlsRqLF5LatfF/YX999/QUBhFcuuWB
b0IXxrWqlC9eU4m1IwF9dQu9XBYTV8Io+vaB3ri9za6OoaHwauuhTi+TIwObtMtfAuxGDKRP6siS
3F26TM14SZIpo6d/ILIsJREIC+y1ehpAIw6tS9L9Ow60h3TIZM+CCjeoYWnW09uO0kSNU0sgPElO
7KkJx34Dfkc2pki9r1+bXKA1QG8kchWsOuopgvoH99az4FSZFtf7qlUagEfFKvy6x+lpWVQMNUAv
/f2U3e5rRWVfPmwt7gRzuGYewh6SX/amvEdKbf9YK3YMa0HTEWQiZ5/AHo28+jkOD5ktFEMa8lsy
85qPS6DaOF1VfGCLbU8fcmM/85tQKu+khVtgIaZ4mH+UCCRCryh1J8S/bkjx2Y1e8ATZn6P+i5vF
5HtAf1x2T+eAOQI0Vbw4RKvOetP1957oXmwCIz/RQmT34qgyxWPRd59er7CKSGYs7Stv/Mww2sR3
5wyTGeftmkfWIPmicfqsIyX4HYb3pzS5exe+ddZkz+tC1pa2UEF+vsdaWef7D56oU+yWdVkTkbPo
kpin80gOVugUKjIa3npYsUlgsocgjl8EIN0Y7IOj6giB5EfsfK0RFnifqk7KV9NenwY9zgi4TQDY
k2GCMC6RmJFEVoSIcTpju0XWfpYMwW/OjCS+p5z/J6UWEVN3NIqiUjp4J3bvfer2AKyuXgZWq2xM
08xyytXgDJSDrzRI4GRETeHJyiUHqsNZBJinyzdCg7or5hDnBD/TnqW/49TuFhdI7VNHhAg/e9MB
Do19h0/0AX7UXfboDRgnnBTF5XZzBWdWabSa9glkWJX+fu4c2+Q43+OD1VCjIPTYMcsnBhpKuD7z
StGLMPVYO8yA5Xj6bi/ocvW+jgy5UvRjzRs3B7jVDPXk4OVaZnJ39M4F7tWW/sUYPog/c/ED+84R
/0ZEaySevltxDlkNgQM73IBq4IB3DAOunVTWonLfCjFwC9/wNRdrB2bQTgX9AKYs/U2X646ltcwQ
oMfz8IO7l0DAHDYCBBJYUFzZdZSQ3+WNLS+e96gxU8d7nX08LuRTgVF8vIhVD3gDhtQZoAqy/tsK
uTRGDZPbkRvQiEMjtGNnOZRo6Dv82lf1VahlwUajvuKn3WeNY3XBFZU7hYbAOUTtv/I1EPdp07P6
PQq4MqKvZEUNpUBwvRCU7FN+sd9tggv6/SjfPMZJqFljTNRzjZ28ft6lu3OQd1KI2rTgTg6D4V2S
cogxIYuiisIWbOS/mHk46yMgNQH5qzthjuAuLVbccTjjXyh+mcGnJVaXJHXipPoyMJ0PotxJP/eJ
NI7qT7PFwFepV0BaqBMGSkuuaZ+YdW2ilZdQemR37GP5244tIcQojJwpsMKRSxVZIWvxcBB5woKj
3xoxy7SaT9uUV1N29/OOJWYHi4v3n38PAlXa3148nEkSGmcKFw+7KrG9xPETezCduTycudbfJDI3
51Pz4JhwcBtqWI2Fn57YeBfVhAnJYwsIcZ+qedv9YDjfu7gMmc8G8TLrlUwYRmUU/IaKCH07Vtoi
P/pMbDcqxAzGKDqUThmuQfcKJI2Hwhmys1Xtb1KrndFqU0Wq4w/SsJOqTxc7QHCCIfMTmReMfUHS
te9g425Yyuo8GA+GseuH8gwL2TUz52lG25Nhp4SB4jDsLYsnJRchaFD7f355DzIKemoo59+AqxC5
Avn0CNmeKvdoVtXwzZyTua3GHetQQULXMNB16HEluyZuW/OgGnJb2C0didbjMS4EwQIuhzfHJxfa
SEQhxIlntA0JhQ3nJEbymx4XEYL4GwFhYHu26KFjbISKRZgDmMAz/5Deh0KWboKaWvLP2cKWn0E2
BZF2nFvrKc3Y9hYwNW+Cf83CpP8R+tWJCXUaL5TAM4VdhXY8mbuMYDfj4UaSGEsBp1iPd2qhtJ+a
tWSZylfkivVDwXF8qqMXLS41OGDOqYF+l7jO2Q6JQZFMcDgzTxLKSsx/9+PlNC99rq+GZ88vptXa
8H+0z4D1Yd8TEczvMCisk89sLBhEv3rM9/TdXQqs5Biq6tO22sD3JN5tBPC5SHzUmotFyTM9o3L8
T85WgAS6lfUg4ZMPwG2KdmF8arTsTUqW7PEanljRIShCI+iYq+mysl1ZR9demwEF2aqrFBakrL0z
wdSP6BPH3nD7mp6JC8MIaZdt+Z9g8KTlLp+aIB6opdnrE+EBePM9uyR+E89YzNM/34M+2GNrHpRr
QyGENsbVCdVeAGPY7xim78X5ymrEDB5buUia8zox/MhRSOVTubQ93fqy2xVP9+JFfNRZU3X4a8E+
wSTGqK3EKLptGYOxeAL0Aodu2HBqEy8iVS5OLqx/HoHOicg9Yvzl7QZliq3nhp8XHL5HeeBMjyOW
iscgMhsiO3dh5CUz4YPNV3ZrH3nDLtqKV/v0xZJri4Faw687XFYDSnclMEFlKdNTuGToxBKczq5v
k+/PhmovxLrgbujNOHVSpYgfia5o6icKl9mCiOKSAkcquwd4uUpHLK4aKyYuroqMkdjkYWuxCjiK
oJedABNyaIRz7lzLBfB0IJC4e5VlXnRm72FMWE1veBo+HaUpU5K7Bwzxo5YcX0es4vr5s/eoaSkz
TncEd9TQBVhx+Ap1Q/xsp6Cbn4ipfpAPTOVQMrZ2FDDxC3nx4HzHE6xE0pLuIwA5BNkHZIqWC7cB
rK1s5JEn9ocfb2bJqcM+AA3QAL3ceXtfHedMPGBXf8WpJsiQyRahRP4uGKOLOXv98jBP2J2WMeLM
WmSqxnbQ9N0NtFgSupkvvD+rCpLmCnK/Kpy9G53lUukqtmxCfEW60/8uO4AwR8rqCs7t33M+CWGm
iBVJpX+7qxa6cvA0r/7Zr6/wrsM+oOdBxmLLkqAhKUDG1u1BjYt+lXBwLVajxan3KsoHvx6YZrRP
X1IVKfBpoSmOR/O8Odf33zEPVUmXSUjC++dPh4T8F6y6MaGLe6yeUtVpreTqB9/1FP4vF9qNbMpr
FqpdOTucHVGMDH+h9REmQQih46hqK2Rd0ap/qlC/+/+XcWiUbzm08LURUF3AFntZtJ9EHIkMte0/
AZaUQUNMikYQ5oerUPvKHGMtaMnJhq0A9pgIH7RXTC1FLpKvWKRF/4Xo0l/yy97Dk2pltMWezjIO
vBzCVPSZqf2v9I6P0FJX/Zk9Mas+0g1SssqfOKL5GEuJBiCyJCDvqAm96POHZm6kxqmY1RVZd9BG
yoSZXw7yp/0O+uH6xJqWEMeDdtQbvPTvZ+jucQnVviFy5/audsVxfX88lEo4GsHc3HG5glydgwFd
DYz55APs4ZBL2wZ74/JYqBwAIN5jx7/z7x3I2IJu+RXRSRppYSpJkHNld8GteVRLYMbOT1eEYw+h
EA8QSIF2q2DNhsm9im05lFFi/m4mqAhEYCLbJrq9k2hYVsfP8d+jqoIyHiqhWWYMyx535hrIDJyp
mirnX1LVJibie1cPETEmJkaBuVG81b2Pl4KEzEA2EQCaJpNwJPfcavgniyN1q44XdXmFULcA1JhM
sO+SiwL/0c20QP6NlEA0tdx3V60OpmUBvjzul2nvqz3zBWVljla43WlnsVypEnSojwkghyZs+Mpc
tRv7pBNJAmnEby6MTywsXMhdYvhDN2htmRdrbaG2vujtxW65Q1tmmrq7zDVL5z6I6Lza2XeDsQij
I8CmUJPNP7huuNbrVfDDmHjgl+3ZRtSAG/VGEO+cS93y7mrsEJFH2bB0nlMjlouwpjmkeM2QwTwY
SuBMh9iG2UIIwA9a57GrB77aHG4zlDZL0IJ8iwN/BYWcHL0itQ1ieTcDsBKc7YX+VE0B1OnM1cZ1
rZ5Dg2bA4UpsDhwIGR0PzQHr7VpLc+bkMG+nrSeHGj8jPe4l9nEQl+HehF3S4yeXN64x1Y7AyCTb
3ykwqJTG2GvfM3rghKMbTjLrm/lb+t/7siSIOLncCy0px4SsJsoh6ExMQs3CoxwJMdsBpFFEhNMr
Lk0T7GVJ+EtrQaZuT5OEBL6fT39qMxRl0hCbQTdYOnVpjhRgmPGAB2EDfvQIsQauiS/HqZYg916c
YXM+osjpGXvtzLcRfDPMj3ncFS3c0gMBXKSSMUMDE4qVMD/hT4BQHI31jABuoQQD3AlQpfK2Tdfa
L3nzcgJRjK/wbpyCKHAb6DylDlkOzIi3Z3Cu+TNW7tN8xSGq9wMtjm32Y820FYoqXZuoUkPOc2lu
YEk8e7gpc1kjFkuLpsnW9gCK8/+3+DhmbDmUkNKVu+HxJ7cqaEcni6YRJSJXzjpK/IZu164SH/4a
UfGIAmJu6p0LDKLxdP3Yp858zj8rWyWIqU22xRcVaiK80JZ2alLeSvyXlJxHD4rzbVmRmZAT83vS
ndLJQ0B+xEkmU7rckqyJdofBSQE1YrdZ7pKnle1V7hzTL3UkugjBtzgfeXelphFVX8mQBaZj/Mmk
FC64g26f8HZisRqgeudBzOq+o6r/SMw23DpZpcR/MBmfpIVqgd+DoCxTI6ePd6rV/4wtDCfyBN7w
wCC1I+rtoR47Y/psexi8v8UsCaaq15xRKky5CAPIhs9i2cvCZbmI5pMehrboamRe5urXFJs+nIye
jLKo1d2GepZu3iEBE4Kfmg1GU9prQ8xaFg9Mrb0X/gyzjAd7bhuSHK0Yp2ODlc47y6GbO0vgb3qW
WScscYPjuDqfgHrI6P1CAHz6yujl4xUAh3ulVeCHEiHf4eJ7LQ8f1DZPZs5ojToxmWgbzumV1+7A
wtujPcflKWiBwQsmyg5dlSMj7N9ttW56HyjXsgNn0vCWrE0AYEdjpTJGVpRHyFdSzQfesXHsrIrp
tNxe0wfWYkkcGDEmp/fNwGlzr0kqyIRVstSJDl2WRdVzHBSUH7+jfnsmvHVX+g9VdaoJ2qNqLwXn
RG4ur1o5cOd1Soq3FZcXan0d6ELx2TtyZx6MBRI5qlbWtcWtVC0anLhaR+KwnQ+dNrryEeV9FMVb
CU6Ohy1SPVhBXFlRF1Gjy7YuTuWpBkAKG1VNFL+G/WeCzUkLu/XRwRr50i1620bGFhw42k+W2lqM
+UMFY8I/Gm4iyR/OY4KsXUx5fCf4m7CVn9pcLjOjB6oOSmgDXYkUJnpjCquGlAoG08FxvLaFDq6/
c7UWpIRhmWki3s9OP0XjvZ1FXzcKhPAiqVyYN+1af1Wzzx26G2iW3vFwPFLVVxO3Vbg1ThYZdFxI
igFfMKYIPU+1ZbTu3O+7m2zps7uTGxBZIEJdLF12vktpriJfY0eDsGvSXXp/O3QC0w84FLbMQYAK
ZzMsTENZ+SmVcjdBUMDmLhvH7w8LULDTHSkBiHzHB5mdAxZD9wk4fdc5gZEUwXlsLpLOnLnnAJPj
MLPZCEMJEH4PpEH9G5w1UNfg24CyK2iGqrh9RsYBxTU88yDzt7nYT0j9FNTi/mRem3DUlfUm13pr
Vx/IYEbKEgNsZezBJqcXLTWq304TCgNm2WXm0766IB90rmpHG46x7Pk6yhCWA/OQZ+j2qrFDBSej
2ITgLMVQD3y329y+llv4zMPvBeIoBcDZBvpYuMeXxYHYMwFU11IzyksefNzO7tv+kqb+q/4npEa6
odXXcLhSaAQap5/GbKezTuNlSb7glR99DudNjagA4jwgPTPT0W9YX+9BbbYGxuB+hbCy2C8WMamw
Cbhd8FmOhvYshRv15hUOzekKeSakPJjEfTa8dULqgr+IT0QQHPtT6YkGJ9iy67ju/Mc3qmAyoLsd
H56YzKKoRBn66ArEBBkFkds9RlWDOY68aDaPS2R6oMCbnDeTLGC7fa12VJ35R9P71xjoa/t/MRSn
l/Z5OniOpNv66FGeR3RgG+71ZDZ5tP/9IqecnXWHqamphbrMNCjc7p5pHJelj+T8mobX65kQEU/E
hpz0F4hKs5hDxm4yRDN4i5X2a16KO1dRmpz56CkAod9uDu5xyxumUWBz+8rCz5Ov1ZMliM9DyZgo
unRY6ZR+0Ac9I/0NlDoOdiHBukYbcrojDE9eR0zLTG5htqAC5m1lQnE2RsaLLaDVj3wMk2XH4Ird
V/yHi4MGlkoVQt4x1KivnstUzNzbHP7sVNByi4d6tIYNQ/GlQ5WMhJXJiio18Puq6a+cyVyKieZT
cRr7BYpZ+PJAwViGN4/Me/WMtMxLIM8J/bYB79ukgwbj2V0Uk/Kj9E2VhfY/q8XA04EhoRprOAwq
xf9FU3xQZop+bAmzQeBtEHNGDkwaGvVdwuNKN2eXaILOShFAnOq9Oqef3ad2HpYV4G7tm0RPR5xc
zEfEHyWoJJJoHCgcoGePcThHPP5xWFajMKonlkpKYM2ZiaH1tqp/bkQQT/Hk5o3Y7Pri/0GcUg+Y
H1rYeO5DROKFtY3+MBVN2GxT8OdIKKZZdeGOD4N1KMatYt6gHjqkb9Gojr7e/FOgyfAJ0+b6pQyK
sq3da/wrioo+IuB5UxEq3sSLCFCd0T/2xHjf+ianOdNcfidAmMYU2HzcmrXQB5Dps7kdd5bBbif0
h8DmZ5j2iyv0L1nr0+QPREfNMydhWRtGElE5kHhIVMs/Jz1f90kzx2YnNjlixOKEEUKkHTkj1l/U
+ZysyVQvpnqE+fwyTf2/Db4K3GFNFOGW405eGuoI+eG4ipFtPskwd3gk4TVLCOm2kcXme8SaCvID
RzcRvUEp8o8G5j9a11+9em74A7IfEBN5gRtVEUdG/y8p3c8x/AAMcXxetX6dUA0mKgvXUY+OV4lT
J/G7fOceq6i0G6JfCsJU4UhkgWNT/KpidZbJyfWvpXtDdY9EXEY9+Xz6ZAhrPTQ/Kq4bUG3ya+KT
iVVJ2np9AJwXl8Z2fM3HjReBJoMVH3SIlnLq+hOhyTVsmOxyejrASqpvPkV0GwjxwlAv9/PNk4kE
puXxBxIqC1MJFzcH4T20jEnIW6heg/LRViDA0roMbWvhq+QB3vb+WlYadEjcSwO+wlf1RErYGS2k
tp8N8Eqdvf/vUU9d0WOzY3YdA93cbgob3iAcKRyNZQ//vq5TCie/FM8VOdr4Gff5md5wLUpvPMId
HjGddpEXlTgR44+LuscM//QxOotvMDUxQ6nj4SY/6VXL1mzV1fPZJH8vxw9+3dtHLrN6sf19JrhZ
yY+tf1jyyW62uHja9BwZtFl7A/pMrViFWsfnDXvyJB2MsUYQXXmuShLplf2P7EZGUQDnltdDHtXT
7GdIr2MLCwxZW0Jwc+R91aDjccInJqB+1+3d26v5bXjzy8f/TmAwqKPl7zNQisyK+nrg7ku36cAa
chVO6YSgxT7wegmwVlu6+pDd6kM6Ea5hTMN0z3rIsM2fuumft+Eqw8Xufv0EXojmYwstWs1cLOIb
Jb7XAw7ApXnF5N7cU2IC/Q8UtR8HjVLhe0ONlsaoaxlzC0wGTsJTj0nHCt7BvC2g4tqBdukqDIBm
FtB266fVOdGArAqNkKx2O5W/o7CfrGCM3GtQhK3S0ehhFMx4Ldpwe3RMGDmMZTJ+uWIEcGmaJFRg
5R/Gu44wG5mXRSEJfNQRUpdTYTRqJXpCAgkUZ8Q6wZ07C9RPWV076wg82YUUgJPXJBuY1gwml0Yq
K5AjAueCUv41K/QSVVp0lF1v8ttrz1EHGGo3vfd1hOuGnLq0c3UkS7KvdfD+5JdimbBc+brrzNme
J8Pa078INmoVXdKlv7Ici6gh3I5E0TZf0/ixTJH/639SobO6djQV02WA93+ZW69xgKlNPQ5T1YEb
5obvzHJC+iAtfAG3iSmf2d86eitGqLLfoARWsNXl116J71vWy5P0AepmAugu7h7wycXJ61G8uDbO
GDIBNQK1FnqvWD2dLY8FnGpPM+fCNHmslM8+JvUYZpRXq3jCwNyvtl1TVK1/MF3BBm7x53moFQSq
YEaAt7lp5Xuwp81no2EiKpzudsZAQJItfPrcgAsm1jfsUc2S+5of+2b07c2fS3X/rVtPlqjTnY/v
j3P3lTWB/k1Ks60RcOEZISg0KHS/RcxJ5FMOWRwDyKyIzOV4FdWzWb/2EiS2vPbZ6aLvY/O886Av
zRSLi6dOEYwGjI7HgbHsyT6KiRQkUBGV1PI6Kt6RY3QiK6lr6z4IKkMXIEYNkpniEHoBDbo1/gkP
JjZ9CVP5qrMG1C9IA8DIu3edKxQ5+vbFrZ/D5RmPOLo8Et7/V2PYabGnl5mUTRRIdwho6XUBdqYd
EupTD4sNQjR8d1EArgJnCmmeHrP2Oq+mT3OUfcXukd8Lbx7nCnxHqdV3Osn+r8QHIb8+9QHYvexU
V+bRB/o8elzh1EbPSWGo4OyfnWYjXmtRaxLlt8fNREEbyDb1MkyKwtox8ZGWl1tQICand6PCgI8g
SHZJ6dvURVYRbbhikxMn2xXS3lFDfiacXKar5eKpWqhzKvPK+halJUU0v5DzyDE42KFqqjtgy8HK
MPKCbUcA26MZUk28nvQZvmol8oITmhMYVk1Oc0OV0UV8ob5MOjT9oh/rPkm6VLlPMqyDlT8fzBQ1
nLsf+IRtqxfyYTsKACUnvWSOtS5ixivUqo5OS5hmKsfXy4hCCEPqqZtCokVhdu6qO4ZmuCCWnv/Y
3zcXHwazZvp6Vl6tlWpsSh8/ID4JOq5MwJkNzltWrwSgGkpIQbY9Fbov8nGAkN0jmQ/AL6EoRN6V
b4ZVPWGhwYH8GVI9voOG94fBRV+aD5ze3Wab0cuJAhC3MZyWfTKvQFU5+gSY1cOIb7TkL/JIXZ4I
BJfQdF962tGW9CBMvkJNDxTj8UfV8vac+C+MAqTtH8jxPMTVS8xBUbsGd1DTPOShejn6QAyi3R2/
mbZo6Vu2cAd8dTUFAXqkTWXibcLfWT/bAqvoYdBOBDSZGP0yhIuBE6t34R0AsAIqUrz0PbdpqtH4
BSSfiB+yRXEZrUUscG/l5+Kpe/dM9eQ3YxFeWKEZgQrE0jWZYrp5oD7lwMD1C5tFLn66LBOECnE6
hlpZFi9euH5cgHeV60j6IPjsRqG36ybkNu62paoyFotiihqnjYpRUotAEdT9OMoJuLNpEFipOm4y
RtUUHTP34vuDVGFJrgrdKwZlgw1rGbinPl8m5VYlPMXyWgVZ/2ey/jEiwJEQ4nRXShmxYUIBZwq+
n/z1JJRTb1FdH194wEQ+qb8X0TtTjaVBHVlWvayHFKutZLiPbuMqox8B8qtWa3AHSnoGMN3SZTr+
UNTcMHqJuEE7uyJncJdUctUj7y6/zDLzOoo+VS0H97n73Hlse2QzVS+6pSWUHfUtYY9179y/ZGsj
NI0nmE7x1EKV7UwX5Dv0vSTSk0A+WqXI96uW13s4cmbu+93SYW/96Ia3zI9qamSyEgD1zLbFlisi
tskM1clzalQpRqatZPGu3wv7IxWTthfz/6xMuxtQQeApROTujNlwYyBos2T3bW8eYCGUPj1EWqHO
xv/VuHK+nmfpMxVgi8fZ9rwcEbRmDpJxIuxR2usihmb1PzKa+SCYYWmamjChyBDSf8xTBFIsP4hG
ZUgAqxLVjKp3XnxWD/aunmXelx/rnUyVge8vAnB4bGnNmd9Q06pUxBMIlMhfIXmXntsJhJ/ZIGgM
sIDn/MR6VgnUxO9GoHx9xcU1xTorcxmMZRxu9ugqul4i3tgcI8nh24HkvkqFEQDk3vmo0JrmQfO+
mxv5aezMkFKMURD6BhkQ1Y1anowAYn2i1R24b8ZXx3w8v03RAb7pWdgP8Ibw22bp9y3ICpGk/FtS
MyAaYuTczK4kzyRfMflOT9Bclu0cY/iTMyuL+zZxYQEWW8XkQW6OvSpiepSacFLO9bKpOudtWgYT
GLSm3NJX3PLz4KEG30HCV2+kZ3ZttKlrowDuHd47oP6M5XkcaB0H8yMlBRWWDKMZ36gZ4SAjYvNw
PKUoT/8XhUXDkRIW1BssLWMkvF659+kcpXBeW33s1E0RlsPbzhK6ZUk0f8RKJxbP2ZyjGV/InhsV
PEzPg9QJoDd0MUGd5ARmr3nmgFjDSdLYgIJ1+0VTzk0uUomiC9a6J2buCYb8IUDX9HzJDrmFxEmN
wkI7pgOYLNQZDdTuqOagHMCEL90i8pYkDKM3/y75UvWgUgTCMtnUpqVjpvKoSPdFVzNcuFWYBSxH
8nm/FmyOQtwJarDkVXG7z4/vntKZFKE0wwJM/WNW/7icurn3ujk5+4ubqldUwtmd24k+aE2wN7iL
YV1P2TuMBpzv88o4nWNDl58mNcEu0kt/5+G6lCKp3LGPrbPNAGToCICSRm8PnkjEk7nc0pPOmXVZ
YB7HCZS9lhYJfSGNJgRu/EF8jQNBqpRObSkV0ac6ZZNHfu1cF7DcHVyf2UIjyg9YG/juyzB8gPEX
X20fUegaYHEujiAZhUmYJe6XZ0AF/hm++d3FwOuf5pAP/ohZdYAdlAsPcLZLD9RkUZoxbHhUjYtW
4IgiJATmygpmx1iayJ5yUqfNu/tmORyfqpCQQPv49RUborHmOMJODhtuaYkT/Iy9lgJXT0EAAMdf
AWT/qjPN2AWlhqsefRrkg+jyYZB8y6qdznjBC95Co1vYoHdvx8G2DSTqCE7c/IrrZGDHnVRz+8FZ
I98LniCUcJSAiuY+LHazDlyXTjM4Pe5lY2fkDKKfoknzp0OeBc8PYSG/qq2lI8NG+SZr2Ip9jYJd
qBn9ye7j+/yXfwzxnZoqr1xAQ4VrRh/O7pVk8t+thyNa45Sc/nvBnXDzOaKFpHNursqpOyM7Nnz7
iDV9aBDgCy7p57i6hlMlhIEEiLGgx5k74GT6EKwH+75d6p1Vj9FSv3nBCb7YtyE1toRdj9nvS0Qa
U+0YRgtZ3P7aAGZWvDdtIRaYKte4cpAGXvDF8VFVVRMGBmtPoQhFRqFS6m+L2W/FBShmf+zfzQlo
zGODMusqFSXiKLT0hVkodqN6gIEVrV98mMyvM4pHiRWcVgh1MNVAkvWoU9uX0PBxXYWhIALUdmys
WNPr3+3LoPKu2zpTPdyq1ozcyIjH1fW9uv+7PM98tRvj0j6k1ZpTsB5XdbcKDJImLZqgFv+LMSV5
7eQwBBzjLwc84/gukinBrHxKCmCHNOpMIEgVjPM8ArwwAGxjX17T6nzsrUSxX3Wn4HzEIV1tv/GV
2qknUGJ5cqsvoG6yJ68GwBCMfrrZvnOM/e3wMEXA/QTwYo1ybdTU8YMxpWF0nkvITqUh7RRDV2ye
+bBAAroV9n+MdzYPLyZ3Q8hFTVkn4ogGnqUAee5XJx8ubHncdPSKd+xw2du3yDxdFfB2SZ8CB9/0
fmUYj54zdNyvHDoa5fNtFxlxr/b69Wh1JxIwpuNZRfFwb+4z12J4Z6CvWgtv1fnWMXwye5ckc3P/
LECAY1W2PLzbfkAYN9UTooSuUNkXYDx1+XjK6aA9ydj37f3EfP2RjqOxpGBJV97JQXJIYh8QLbDM
LaZnEgQQ0uPuW8X32FRs7T7WBsxF4KIS5tTJbgTKyQhPKQ/b7m2Blj8KEz/+H80MTVfNQL9MfrkU
SrcGExeov08XKqrGiEDhyCFjCy0caLK1S6DtOCagI3vGORHF3TY5ZPndQAe4c5TS2xfh8KDPkor7
r/F3EsfvBS2z3b65L7CD0QZUhEaIF4h0ict4JrgpnvY70lq6Pxdz4dmB6pqyzvB6xjbEFShyr+0u
gI1tSmdB/Pp3h3S2+ogIqbl7gAOsDvD7Jvah0FGaMBT/w3CDMinxEdMnz/8ROYCf6h/5MrUFVkOD
LksnTZIOYY4mCIsVnXkOEAoRqnlQslerPy9yyxcxjkPf/Ciw0TX4Ov812sR/rWu4smVCjpzHJx7Y
+a6DeiDTxXitNVX1o3uwqIYXabcIuBuYOpZDow++OwmPcIbadLI5UmLjGVJ5bc5kve7Vt1MbXdzS
mrKe9AoXRA0bP3ne02SJBUCEa79FCE6NV2B4vgisG+9A18J2Ci+oK1Jc+kjYeGqsZCJF52U15yXs
YW1jSS9SydS/PFYqcdKfotevgYeZ0+51JSzDIhYLZy8XlCcbnEl3Sa7uUvQYAxn6V/NNPbHMt9bI
2o98E4LZBMNjdJiFhzMP/LTrImlTHp2Ia+e+6C1XLDmQ1N27lrsqTvdcI/kFt2pMZkBtDtQ77cxA
NHSBk+gMOOtdDJzhEfrOtOGQOdlTlZ6pMV8SXb48mgfeNaSxedWALHjPQ9Z27501/Jotjj43qJt0
VxjD/6S9KL5ZJAY9XcU+O7SeHwbLme8JjN5+qZ853zogssL5GTDFSKCKnE3Xfc8qyFxOa+PHlztN
Q1OYbdj37VsF+6IJzo8UTcv3eClU1S2vnP/qxCukpM8z805pz6xNh3qkK14upS6rZqfHAxZfbpyU
gKahhrDIPT8ioqEaaCW6niie1tdtk3N4jviiw1eHSMkYH/uW2JdCyvGVR+EpZf1Qux5Zzh/rtE3U
KTWWWtyY7A+YXtJQserWJaRq4XVaQyS9umNA/Kd0D5f2I9aSKXii48yy/zjrYymRCexp17LL49Sg
RXhFpWf8voCGcB2Yl5HOJeAKK6Gjh+uTPwgZuhjdvB9iKhCsCqT9inSiChlvgVcOH/cojvv1LjOL
t6IO+fAxjXz2z3mAM7mGDPfQQRc5jvqdDwm5RpuY2dbN7cRuAyjc9btAdsby1cn6dpMc2e3q5cQJ
af7lpI6zXcsvCjwWOwGcEVapsqzYNFO3JNcVKHcRer/UiP++COPsC+r+pFZlGXLBJa5WmS2gAgoL
ZgktvlzdxM3Wful+V/ix+Wj5ZF2+D5X1lJweOwborPSmeaAWr6hmt6oJyoN2KWkezR4XunVttJO9
Yn2LHxlYOlpjLrCM8MTVZ4RNJqazrKtn0zb+r9lBqGhczR4WyU5I22lL/TiTvjFvQ1YVQ42wAQhL
XjrDvC1jJGXteY+7eo9e2Ga2lfQ5C9Hjc+oqEPy6k4GJFrxTH5B0uinxMqzRODIdO40YnOoMAUq/
XMjr+Lp59qSb4xU8rPeNCNDU2VX91p1s/HA9JgATm/xhZ1Fnh/HhnHEjKDRR2+AJQHyRp9Wb1Q14
/LMMEonVzWX7Z+NpNqwBGM/Tx5GDUtKlg44JWiz0NwXEvxZe64OR+1i5dOPFNoPJrQmfttq/FwBt
FLRrKMIL2I+KN4onPFSbIZZbDxn8nYnytMfHNMIg06KMeZGbdVvLrcu+QxG+jEG6ZiZYmmBA5usb
8UJ5JXtuhwDnoI6XMJL5tJukgjESkRqx655HhwtycmzYHie52YtJJ+VJM86BP1YsBBpVdEVfQqqP
lZEpUflPbZDMRIC5W8tFGcGU8fo52RKd+F+eWT/Gd4rSu4EXAlkbtvJv9/RJyoxz08qjceCOwPkM
lhABBdC5w9feKRzOUgry+A5gMcuR4xPgqHBeO1XUTfSJdSfiKFdIqeFZslTYRbxXtPiKogI2veis
3S7iqFQp8yaAIdbinbQr+TVibO/H3PEX9pkX23HmPl2PN9ObBIQVpEko0kmeIPxy0vdglt7fZufp
I3l4LU4Zx4HvZfmFol9w3dso0C+mmgAhbyLREFCGVFGJr4U9GuBzmifUXRcjMBw0llhd56zYkDJT
CcgExBhiLPaV5P4PDRygidr/WopA4Bu9AfQeNc/PdgifYmCDVZgBOSwH+CrvQj0jj/HtWPb5Vxf7
x8OzGncer17NPdvfanSZgWcSa2oeg4AgGCU8cmeDRXsZZtW2vzIFFMPd8bonhY0YTYb9U4rTX776
GttTCbPVgczq0iX9myLDu86d1XwaB3yJeDQAQzXncwZqLHf7HXhLDHKCp8bGf21gaYjk2Nlj3y/P
xTT07CCtBKMBbWKv8C5yzQ0+jFKaKFDjTdjERKY1SvjzoQ67yEn1r5VhVYjh3FxdbXXkwt2WpM0K
NvGhHNh5ZTKCjQcimjggmLtTgUz/paIG/VIKl0qJm8/9HKuQJVJK/mFEe7oITiikldmTISGmqb9b
ze5WOSf5PdPz4yGNYg5dqH6upLRLZ3khANZF6e4GoeotHWjOLU5U45CEJCgi/1+16m742yuUd049
1IdYG0y8+q5b1+oMzy6e0aOn39/98vFrbKCjn4fMVYWwGyyDjrG0PPLIOLopmWLDyAlKPeaZXTxB
yF0saVh3BoehU3H7nWJ00VtEJdfzLVYBiHV3e3g8eKB+HtyEdbrlx5T6/MUqM9A9iPb740mTKQE6
iHXQCY/r6FBDyvalpM6uCIQtsxhG6e5035OhGni2AF1mr9HJ5mctMJ/o5+VvvvoMCXxtz5UgxYQY
9Jrz/kKTEBvI3KEoTz6Y/m8Zct53Uosel9Hkg1jePkDUmG4ZYHYTM4O7WkSaBOinnAVN0B2FlEzd
d/bICpcN6+EtOgrJ/Ibk+l2jZvRWHVJyECQ3M43Ir9mplIloCzJ8e8BkbsI9zd5gaxHZ2YQfcZXk
P2XyAXymaJakOniOKeu7AvHmeHOQrdh8cJh4W7jdc9D5vYSty6c11TQTRuKLhTSd/N1Up2UFpaxg
hz/jGLqyTsAndzijGHBhApLhyXr9EXqCoOKR81MgO/uEe+A7A4kTR4HFxaEL7tBwNN8AiHYP+LJh
aMKYyRUAsY9ml+EEzTHc5mfMsF6zuTfMSPUSq4tDkWyMKrJJybeyOn7DuvYbuFfirLGe9PsC24UR
mnCGz/8w4mmqO6EXHDKkhMs/Pj1qLzI4+b7kS9/l1r+SUCYom4PmPFrVVgmp/G7n9NJNRMLoUdUf
y8olwVS3BCIYk+oiHGsq4uStZkoENnaLES/MEPCV5emOF0lhVj9InYCE79dTHkkeOvwbBDwx4Fv/
5vLLQlGZTfrFOehgD5AU7fWW339CaqTkRCyf0kbN1wscZCFbojMHTWPGGWEQd+/8crYc+yKDH0Xr
f+A2drSQHJQ4o5paFLqb3iegJBZJFZhNxtXvpBhCNjeXD8uVGOPI+TNGPFSO6wIkRSA95sJkuE2D
TTFdTVJbu5ECc77nwro+QBYBLIaZ6NnGXPVCh/bkfJDuXcpxE9ScT8Tk8ZSJxO4z1VP4s/pOQvlY
/AdV53oSDyeZI3Ext1H6Nw6+2B2RvVx+WR54Vtl30jU2HVzfHhoSLcpZYRLrVHU4ngdZ4dWnionr
BCXn3rPDwdM08p7xohZZg+QVnSk88YyfFzMGtKsmUCsSswshhO2PJfXLnubdMEStISGuPpIPTnUI
a8Q4qGg0wz22slsXu/cRAdgyvvMa2nJC3qUE0+D2EVkukEPlt0r05iziFe0VDrbvIxpNZqxrRAMY
FwQkhWheojl0Ab3BerQDSlOpRb85GpXzTEvHU9GEUnDZTi9TToFoiTCWq1eNtguweqsGy89ZSPC6
MSL1ZeGcutH+BuxPzP/M0xdlDO2TT09G8/j/pTRrhbSJTMQE/GYU6H/qFJg5sbhRALI+4cCIu5WR
kdRfr/B9YgrmipqKk2R1HNAmYn2AiVq/uqxBYkZLfUSRErZQfaWoFwyfDg1TDgKn/5KBT2Hp5g3N
hWzaN9P/v1+GJQwOi6KT3iAbGT5gUdn8EdiYQBKa9uGM+V2HAuOI63QUBNLo7Vx1T/bH40+HNW+n
PoKqmISmgwfp45w3jy3sTpOGoRtci0snG1URAS6Zco0TtY1Ep6dYku8KykmfkVFlQO0p54BOatIP
deqIyfGjW29nXMg+dlTe1hwhlOZYOu6rHAMskYp4LzK7EbKH86JM+az9/nBgaAAetqBiZt1je/E8
kazCeh2Scb/7uFiFyW+nlejT+ZecjCpN35UWTU5Jlif1OGX2zKJy48DCcqgLIHbA9pQPcYU6YZFg
HNfl7RCz1Q4sLGiaa1j/UcLL5bHwRTV3lfgZ4LsFm+wEG6Y2ok/qVTWpP9f6Td2kZg8n4IGsBFrx
c6VkWNP6+d3dsMWsXSxgVmakb8NoEjaxh0jZ3etUs/wpkPMADw58QFlNKs0HrQ8uSTtDsyO+A6CH
9Xdc2d99zUmunjoGvBVz4BP5/wZTP4QWwhsTPgWWZTE4oMh+lE5mmMmHGhax5d/qr9GeqcIRp3g0
xQGFdPgt0lS2m4RrUN07sE056K/mwvEaR6unrAuI/r6Y6pPvaeFAnXLrWH3JlhxPWJ/83njwhaAW
IBPISmQDG5YIYV0y3PySiwZJzHgsQ2JBjsAvUs7gR2PmiSmzDNkTX+SwcObsG4xV1AIQ+CFEBPVI
EGNQK1MSDwdCelP8K6onhvza9lBfZAD4LxTQw6UlXtYned+rVrHKwFdmHv9Dspt72o2UepkB6zfM
WTP/kK5fKyIhjeWXpWyTnbs0bJFkwnrFCgX2UDuog4id6jbcOtEvSHMLNUg3H57YWDlFlp/olc3e
BmuEJIKCGCJVl2d/Y9LmhYfyR0KCUhGswaG0iNKxidkP8eefQrYD3gToLKz827oqv8AVcRZdhdgN
kD05r1ONDFAfpdI+EmVNFQE6o+1qtHRhErCPDRmvCTkmADZHuUMwydH4LvGGQACi+xdtW2nrpSWj
Oh3kjhdKYfO+8ophYWKCWNcAK9D6YyM4o9c+sBH+vg8vc7D8I5aGtD6CSXs9bse479GU8NxvFUTg
Fgp+svi5kT4mk/LAIBlUPRT0/tilelYNgMY4WRPN9OHGUhyOp0QfikGjDlovYV4HtuSfdgUwF4oj
A1e6c+ceCP/Oh4R0gZE0BeupmghH4u97EqIyr3Sz7jBHJe0fCM1ETTOC9nswGajDWqkw5VWfpPdN
yeiR0039XUlOeGJkk862Y5VTY04lytcSubXx6UI3E5ZluiCztUn6BpcmILTdlXx8yoJmdxM2dNtn
UUpG9POFLe9EMAhyjasMA7Z5W5/rlZ69pLlqN1N5HGtiSucxgnCJvRq47fE04bmzFUuX5T0fFEUq
Nor08HWSMxdAnfp1NeZB5yfW/39lnJ+3+OLJnyEuMzU+uOKUD4spKKWMk5pz8KaV1yS8Q1Qnvve9
hq/7xbnZfhSQ7gCaFGMK7Rq4J+e3vdsrqZXTUOfXscuIooNhkSeRRclp2nPDK4Tk0+8cQD6Aa2ei
tbcqNraBezl3oPVF/HVrI87wd7PDBUNvgPRB2x8mrRZz9S5DLex4IWlAqIH5DEyWzWmlXUcs9FHn
J0VLhuhRClepKaIvvwyToRmSgyMMHFFWmaLto81bCiiXzCkU06BAYVP+3HndTyjNdGg4ZETeKmC+
HZ8pWpt3h0V6aa0CWH+NU1nD5UjYmnQ+9CBj13bwyY/8kSKuBhwtl8JKAnx/pWSo4+Nhk9IBVKlW
4QxclbtFOV3YbWiolu9vZeQrgB7cugwsgS8aGbSLBz0OEniRMqedQgj08Ro0K3PNNjGqI/lwpnIn
UrbYLCoTXjFR0HffwWAZAi8TbTZ0+lUYAEnU5bfGUyb2d0aWo/Dd5yjnFvrf5WCQA0jR9lK5u1UC
Ln4Aj3NCjcVVNRaifEmCwezHSOZ87JlJlM6Jw41C3a1DaIfiDrLlpOiReKANCmeRV24Nvv8xsgQT
YJneZJGctwDe1gtjcbMpG91lNgA6pL3oXTPxTZdfm416KKPzgQ8u+2OGS5JGyeeO5aH0GF7+Xxpb
WMr3ADkQLqnGPrxcRldbgz3BhgMfUZih5Fo0Rstr3pZr3EekhRkSYrh9OUTIprTLB79jdYNyLBfm
2ap4cKhed8YITxPDBjLiCE5oN8LFQ2JfzacZVJbJ0L0ojLPRykuBBuifFWc6i5FkYwNLpmdtw3r3
49pSfLOQ6GFNeXx3ulUEu+s/KW1WdCBBpD9xRfbdv5OOCGosUb6LBEydm4WuIcrG/ib9O6SecK/H
0jHfUESZ7AN7P0ETbRMiQlSNozd0FLG7cHNu0Y0U7Rh74bjDERQ1izRZjEaUM1fnIkAAMGXlDbOj
7oeQWgunIDYU9cCM9cZkaCbzkY8qw3R4jV+dVuFro1RzmxoubsgQSDg5NSdbLnMHGJknKdBrA9z/
IaiKZGgkQLbXAny89siQs5WLN9VvWmvolPcwn0ZRLVlOmZEernTbszS9k/O17ldaNJsXMvE0Q4k1
acpdYQJoTHw8fwxscew4Nyrr/v2+oaK/FPLGg6i2o+gYOf+ifpvmGd/Lu4PLGeEQNm/fJBig1dn4
7DiVz3tUWUCY5tAJRn3IiRDdYWzR6Ze5Qg3oXEVR++mgg+Qzpm7M1oUm+JYdXtbYHIYnkcdU7IR7
9ZkCn7HXPYwWCf8bEx1lk8R302Bh/69XAo1/ZAzzB97dFoR14zmGl+siy/oAGlk01xGeavD3S1si
pHzk0CF4bGFFF1DN6F2X6Ufr7JlAPEFAIGGD9QsTZGZqfKVji8k5BLUL9sxp/hD0hcE3GxzwqywD
E/vIC/4sFvCNLWbbQojySlVyeugBYktEW0xCXdZ6yeK3Dn1keqRyPKS0/CnjkLecgSBwrgNapB71
VBWVTg9K2hhEZl6hh2lAvGfILqtFI0uWw2LioCYeHL2SzqO+UesY/XbDJIa0zXZcD/ykDJrvrJno
RcofJxGp9S72avZX3H5o5vlnssDCYGLyuqPltGl99MRfme5JTqB84n+6l0YcZcSP03fqWMKAJx/q
Jul3+rvNRMejJPzAQk62EbH/xVwNr1NwfWkCk4b41zQWsOxoBfZ+5U6MQvXazAZIrbcaWOtr/QF6
RiyGoeKjnvw1vjUYS6J6cPSjc+ukIA8d9p0cJ+Ykdd0uK/4PZTbKhPCM5B05UEmCdAVQuCheKRF6
rOm7157ti7u/DfseH/kU/gU7nHsZzjJH+ppNKUVIeTdgtOoLpGJpsEjIIkhRbHyWXv/lkhYNnc2S
SDczwOFPzz48WT5db/yOJzyKxmAfxspqT+wmOsiv92Jg74fG0keanJopKH96vLEhkVino5fDQdbO
vgu1tEbSoO2KeqHUGAPeJP9r+k0aH/IyWOMogqMfOWm+DqY8+q+F+i/bBZRufBiWpEXX7IobLdfp
HRP2pOPm0kWbBWbz1RQqgWKa7Xaz49U8oy3UIHgKQ0HoupULY9PykV1ynoV/3PXxDhM7fUNn48H7
uM8cYbZBt5JH5hHtNfV00NPuaBxA4nPq682w45IUo+MgELJ6+MScBk/n3zbL7Tmqb0moKhE9IbOU
Fh2TERIPh1h1NYxyXh9FHsnCJkdBhAKwTzo03sFHiyEcOR8DaBToebMqTtKaQlokz5YvQqQcmSfW
pxQH0SdQbfhvLVAnWqYvKLlLy9e7TkSZd4tAew4V105ZqEuVo6/2NdMuZdb4VCI53CPFZ9xWXxEu
PPd8j2Biz3T633TYEmV0e0NLb8zVxBqTLtko/i+ljKEGPADHveMUOOvudVb4rVBlTe82K58XXge1
QqL43xDyY+C2bmdXBd4X4YnfArMSm8ql4sIXeJZMGwfaQwjizTqL5YlJitVl2Vqt7+eBolZyxXWB
qtX76sLWsdgPiDDltpU/TnR6M/kdkKGcd9EQlzwoHUAL1CXQIBEE7Fkl+7S82eToklNw3rDyCcmr
wqXL0fHc8uAMHpfxvCcfsPPcHz2msh7xAshPv3x0xKDJidMQ2Dcn7eGoHht0xWv4DHWmzQY03Tlu
UMslCcpsCbLo8nEBJ9yI3qkOu7nnco6oqQGbAeb7Q+28mPlpWTQznVyIXfOVxfnODBEXzKfCv6uL
zKMm+/2Ty7ahumaAa/nvnN/cIkP84SaeaQZW6jjUxchi3AmplbU1gJ5SdWR+AgYTTmOEMUTOb49C
p1LOfVw1cVL9T0u2qZNwSaXpvi3A4R5/efJNIXip5vilZynuA688zvgOAA2wJGoDXwweNquwKNb2
YI/KaAGa92iCwvtKNbO/K79/6uBfvn1vvpurLTOn81uD0a5bGGoXllv/LyiI9A1za4R0mSU3hr7C
r4VntO6Y7TBM+aY9YLcU2zc++dSNqniOKAMMHHa8XtFUHFLlYJxr+xa3DWUsnqRjs+VcMahBGM1e
HbVghtKUiPE2DEhvM3TcqYvmQGm1mWHrdOhCooo4FSRO8ArucJQtRgxa9D8Lns516Qlr84oVl1mT
pLpmg4NEnKI1c6uPrpkAoG+5g85q4ZrawjuARksDeMtzkPTq/G+/tnJ5vLALpuk4s5mVbHkc+22o
Dc6NARsDcpkcDTz/1aVGXbxAj38BiyzeoS4m7Ckj8s7TVWJFipeqSb2zny7XuX60d7csuk0Fi+x5
GMgT6Vwqvo7spJsj7lTe22oWnMPJkBLSyemTuw2uDYLXzRf3t9UAJTJz5WQIgHjp0rnAjXJdt/E+
Nj95mYym3FaBEYjQ799rvsZ/HgVktLIMeg3SoTr+qHG95InY6fTzkgXHPx+A7qYIqomWteIz9pgI
F4talFBr125HwbN/wkR5DpjxDtnFsUhQR27Sgw8HHah1T+C2QWz5GFZoij1g5cq6Ookz6aH0WPGe
WUlFRrXA1FxkQEXv5yghG7diiR/9gtSLkhNpHwRz+gMGtmOnYFhxbvC9pwtuUsUx5TFAUQt6WmAH
GlkLMqyE06BHClWEkxJkY1wPFDS/1C3UCRjyCt6NQ3jG4qpp1TDVlax+k5q/lgeXIN6c5Rd4YHME
PHFklWr1RNxyVTNaQJlXI9MHImg0wyvTrIYf8naIOCqtI/5T4bRa6t8HjfiwmVimHsvgoHDAa2rf
bPiBibFmX9Mm6m3hOCSYsPOzGbgxS4wbvRRdrGjxuH0mtOh8x/U4J7m0UkUTtIo1gasvJNxC6B2R
jx9Aj+BJ4Nd8c+9WoFtRC0RACC7Asjm2KO7/kp3w9BkFukZIil2hXdOpfKIMBDMUewxY3Utr1hzo
9j3CZlGK7lDsSdCqeEps1jDfgEkQyvfATT1gFYdVvB2IK/AnpHdtXdQGoUdu9zrrioca5JH+//tf
cGItxwTRmDYHJmuZJtQo4c2CrlUG1WdWw1J3zVOwFFr+a1ReNgkTp1BTTR93QRzZvijzVCLuDpdu
lndOJdArnzAjxQhYE+SD0RQIHXocp2C3NlNkhHICYEg3yBdoFDqagE321pw3Kd1hWeJ+3aHzUTkl
RFcC71ccTvLheXEiD/TTUkXnse6Dmi+/WwYdR8dcU2TaLY320Cz2eZYQQXjXp9NVgudtXrER9TVb
+MGs6Z+RkjUIpjddm3HXhAPhqaIMf8cH/E+Q7w7dTnX/zjExH6QZIdJG28Qvpk+R+nwZKQrWSiOA
UiLaFdQAMnjWzb5+TquRhPwcDak+Qc1tY+fZWm09z+nUc9PXjQpNTygadFyN7SM+MtBN/Fp/qYIS
kxR/GE4uq3Qz8PQtQumC2GfhSbwPymEXjAD1r9BU50yw3K14aoOERE8WCzzwR0+3nTd82f18cdZ+
4bhxBbIXnWRTsh05ZcKVmBLY/jfgnam+jpOM4ZelWgfdpy2eH4cCa8RMIIBG/A1O/DaldphZhmUf
iC6j882drWzRBeR6ady2DwJ7dSDQUMDOO522J0ILX8RzKYFb8x1nGP4qnMEwyFKNUPH0mS88vQxJ
jxzmknXNuO4pW36vPvyq9inev9MGkMbk6eByHb+kc3Lg8lb4BEUldOWOOj/suape68/x/M9XY4Ip
+ndkeIZM2sfIjam80ibuO1nuqvUcUquKLmsSYAUo5Wk20E8fTAWSCmefq8P3D5/SZ9xegVnfZFc/
+ppOhhaJkMieL/wyTL/nwI+ekxXKs6cfGRY2tdT77Oc2plW6fnKs4/RPTTCcsuSm1fC9zPS6vwaG
5SguqHjEcE8PTr5/lckqUNO7kVs1+MjKvvr9ULsnBsxC0f6zU5HGxzcXIJe1O+ZWaOW4VdC7lXiB
IXCMdOogsgbNAUVHPRXzX0Zw3QIGwjzgfC7gKmvf28KeI0PPyx89pTg96wcipMo+kfBQyxVV7QYV
Zrbnq29y/SOwmmZ69KKTImQO3HzA6XQfmvVH9qf1kqbkOOH6KqolAUqEw/CuAb1hzFmgE5tOsrs9
n/qVSIXizO1ecS/xFV23/7S1x693IahejagMYSrOIgFafylRdo6h0k/Hz24l42YOIL4pSmG12WnM
avm9/buuE2p1jgpdbO38E97H4ovrUbeoycCCQTomOj8M8+L2T9b0zJDK1zXyDl/bsFN2x+T6P1ym
yMOXmR6u3FuXTTCwSqzj21aSoAtfjf1HvYWlg27DYw1dlKxYfjiKp36zoSRZzY/HxikhoCSoq3AP
L4MMqV8Tn0kVMmu0WVANwgHjXB4qDqDCjXRUFbLdqOukQMFza8HmcFdxMXT2tk2RuMpbh/+XrKbu
hmE7Pbr/jRXz3ebFi1ueAMEZXMo3Kdc5ICpjEDF8rGaJgBxEoeua0GyB2uq1eR0vDaa/98zJlEIb
FbPvTkBQuPJxsOixE4z6KVIfU18RN7oWsM/Nf4/vlusr/MY1X8T8DtPEETvHXXYCWo5GTq0VyL0e
Wit1VFptbXzOgxZtvI63MOD7+mWzLlv3ZjoUcz0hJ8p7q5unqTi+FCGigkV8e6mREUOh/V4i/t63
ocqRyu3zWgABxBYeQrwsQ+Em4yE/MlUxYtUgtEmgDnEAQq/51sOp9K/dPhxr3GbRSnD3Q0/seSyX
W75u591ZaOOdWYhZRZPV9MdItq63M5xNc4XUUSOb9Fa42cayRpKzBxg2VZO1odSx7+RRmqoH47+X
DIQhaiYWYv5WS/8kluBFRKXPUZtzRL1XgU0QrVtXfE8xwKIdKwP63bjbfTa6bUl2C9ID/p8w4wje
fbUJjvKEs5ND/HnUhynXMG4ihbg52vnljEZdFiASwT20L8w9CCZQOsMRz5xZDSrYmxbqJZSZLeTo
nRDB+zTeRDFSJ79wv4X4lGVQjxUPsNRHm/gn4f9cQm3OKLLN3xMQAus+9LFbNZD/xD//gWPxtI1K
cy/n9x4WOYrPy9l7qOMLurbQhP4LVfdQA6O8JLpXDnuG6G7FF1W43qd315nBl6sYQPvv18O2DMjV
tkggReedteFfJh3BetSmrpZjw5z7+BsHyByNgmjgE5lq4ZXh8AUmU+2e/UGMmRJHJePdROvzIrg6
wEbW5jVWIQ/Q64JBJ5W6/LV4enphUDpx/pcaWq5RqYOXW1ZKuVITWyvYfzzrnI6b0ae76ZZ8BaSZ
0UmbDYTzLqlOo2IrQ+NC8tYWg/lSzGhB29ggfQJTgdCumGZvpfZM8G75nlBV9JjYLGKDGVovEhzI
1dlnwz+wg8hOcvpHAXZcI9O0+xSiavKMfu9ao0rymUOlbrfyvbFOiVKy44OpqeDdlzK5xHBdwjlX
CKKIX54EPwmjP+OTdZvDH+QQSqgZwWEUD9/PLtT8/CJDjxS/lfUExg0iEdrBrwZqbFfTmRBDaThq
qmftwEZHgzRvUybMg1Vs5T0BJNUkixTV5R7EZoHhFbJK6Wa8M1cnG9QsNT35UVQqk4P1VYcTleR5
J3HwhY95ir526TIjT2JHngiEtYtyH5q0Aqt6ZvSKfBp1Ztx9xSQqOABz4PMxMGRX56pnMXh/bTOV
uyGKgZtY4nIrXA7mVJHItxES4hgKNG7MD9lqRksto3PZjBQBffMV0yORQB+VK1nLxQ7FAZQYnYIx
Al5Z3jGBP4YRbE0bwhPaebix6ULRYmANPK/i2wpxKsi4ZPbZIuQwrKC07y27oA+OcCn+KQA2EUND
vQl2iMazfjA/ODgvCZUsgb9K0RlkQxrYNN1QjhTlO/LeVD98CmYjexa3oE68LoMDKWK8lx7QEyXW
Q2VmWkk8Seo+s2EKlWXZeB1G9nxaS37rPEfsh8f/72OgnQ6ajceC3pwv0DbekWodEwhSPCsVSi2+
dTbG1gtxALER0gRZ8mtYEgoiCudqWmm5ByhZlSmAETsMCcTFySZtSywjop2/N4Y6pGNNeWp3rFTJ
IIuAWseqjsRPq1IwRCp+mlMG3FrxKpimV4QcVhS+NSo9Gs40iM4KWl+L/Usfi4Va1Bai8mXxFCcK
i+PsuxggsknL99bEF6dMbouUAmOQwnMs+wdSggx2obhue/ZA1O2Zt5lcBlUjFTqVriraUqSCCujC
aotKyi0bUU/eZ76drX+fzppmIkXrQZoSs+ECVc3M5yVnrwjA7X139dRlXrUqPS/dcITzq0GzHGav
r9Vsbs3XRU1xJq/TXRyDX9Wf6YI0vF8twYm1JpZXgGPKabiMxeFM+bvGV1XV5uOZCxxMldTsBtK1
NXZUWf0uFsZ217U5mVLoCUesYHCkjV1A74v4Xy8QhgtwYmaWAonfsXrBC6YKvKOdnBvKBadD0xgc
DuCCufAyYWnQ0JQeuZDTau8HdH5bSdxHlTpXpLYUylml7Bp2bM/BuyghPdecJWNIVXuDbv2ea4B6
ckYaid36ttNX5/6fxnu35stS6Kr2DShKYGZD6f8t41dzpcAEiDpSv6TeGQdjTyr41SusLNLYTVba
j+jbXoLxHtsuGHvG8DhE1wp6APvQ4uWwQq9OmBQfRoGblHoHhBiH/7gNyCkpWFiUdX8wzcVec+xJ
tk9mjG6G9LDn0fjuk7dkNkhAijAEaCS5yVIyx9n63W0KWIDI1fEFeYO1pLWVIzcD1lzW4jPKT3uw
eX6UMsu1fiOjd1gG0x6OSfMe0SZQbRr/LEAXGRWu23YysW/LNpTnU5fHqfu+TT7RfwKDII2/72e0
njwn1lqW6bnVPYepE1sFiODDwHwWuxd4fTigBxP5lXuZRgmVao+5WGSJWnbLVxsO2+dlDY3Dqprk
7Cvfj3s4q7zIE/VTB/1B87M7Aa9zQwtqeLlZq5Pml9Z9Q1fkwo41vCBLD0/3x0V3GEtuNNqKuXyh
953L6j6fyBOofV9cH3my+IzrJ9IRMR4CXynONsdUijDXT+rRneLFXVOkQs+3cghSUxgWe4byjIWN
6g+/yKhTKqsGU8m5sAbHeRbfa0SfsYf+/oAAY8zuE5QJKWDhy7R9u3FQFvAuNttrcOt070S/2bu4
a2D9QYd/QeAMaHYhmqOMmvxzZtKj/BU/8FIobPzQH3z2tE//qkLZH2ZABwuvxqXgd2jUZ1El6x1w
z6UklYIuvoye+TI4g9EMaSL9v0qfhQA1OzhxYkdBriIZUIk4QDIDGIxyfOuc281pSE+N2XF7MpGF
ym6TkJxibCEKm7dxG3dDnkkuBTi7dONa28T2l32+BG+XDPshWm87N93Lhp8t8untkgdRHke5Z6Iz
mBTTxlAonftcRaYt5prmiTwO92qqmJLFGvi1bVzY4VsoX2CRpUmYwFIXvyv331eXmvO+jMx2R/Wt
TapVA/UM9wqWC4nujRqNOIqPEnllkOqkuggNQiUeDTpy/O672CmIJnd49lhVakuZjuQmKr2dJ/Du
jeXvBKlOaf40gYxwRee95oljor0exgEQsMzxyOui48nb0Jbvh0vhg0oaxsQkpzBnZEdTSLMMOG12
KzFEynd/nvN7W/rGsVkkdQG3lR022+Rl3VCosj0ReLxzRG0r8a3jOGDj567gxUX8q7vubEG98RgH
bXgBW1L4bv5UBPpSZhae7Y6RsmHu78nnPQDjy77aoIqE0u6hsVCn6M9cu3IJ0rs+Ia5cEtmBbKhZ
Uuo1YWKaZIuDAsfm3O6qkE4r41nwwEe8GTxuYYNiR9f0MYtv/1SU4HrNaQvL/mT8BdDFJj906Dv+
6P0nKnTyPJeFpLUx8z8TEy0gqSIKxcY3zLEhaQViZVD7ze8s2++IvXjSn1rw7HSYH87tVV2IgbSc
dxcXq95LjGNl3eKSSq+/3NgKqVzIxr9QM0jGKVFl6wudvVY3gRmt+yMFJuo4zRVckEfG+1jZFnuU
GVskMIDiDjLkfEb6KV7Gejsg9D7lI5iNk6NPwvpdn7qImDel6raMaIAqRnaBByAi4zs033C4HkwR
fLxHR0WkL6H04z9Q25pub5byVznZYEQV4UhiQYJc95zL7+VALfYkmD9BkroEYWHHSaSA5lOs4v90
hxqFTlJXVUEKBWE6dopPkA3dIbJQH09hivFSeYUWvdCQRDMqnkaB/rRXUjspJ1MgK1XqlZ2XDFnb
Yql3HEojbJPUCl4zhyKJyVxUY0VusDpmWeNpHqxvf0WEawHMP9QCxOsPgTnlk1DkgBlK9qP+ojrj
SOiDHHtImWfgJSCrh5vG2pM4ljijs/puZBP9dKac1v6XZA6/vziJh5npFUp1kUGJLodJSma8l01/
/pgHH97y/ghI+git7iiS4qJOg5G+sLDRwO5AulrIQ6ZFKVdqIuQ5G/+5D9Lbl2diKk+7EFos7MzS
EOWDKhnxj+jlbCzSxGmfumBCPmzbpxu6oOkhin7Wyw5Ducty1bGQtMgKSDUhY2l2J+tsO+i93kIq
JKPYTJj26QcTbXFxsjr/eSyjXaqFiFszoHDnnxbwP5NUSdjT6CgxrQ9LEZvb82Ww/vB0k3T3WtQL
vO4kL++osKEGFKroWelL+eO0VYhWifeMC+jR9N2DsY010HUp+zicr1I+YK1W1zKXmadzZgnbGCyl
jnzvGslU8OGSvbFeCXNo6kwinsLgjysz+psObILGPXphsjyRZBO4uigZqlElg7TrMHX0BcxoE68A
Jf4jlOOju/RVSTHu9dxuO3lrjSGj4wmIYKoACDvutr4FYdgzexFfr7dQQN/gzErQnbBZfKtdu+4J
CHYW3uUHiKxnL2ztJ8xmcLaPZWpUtwddF1NfKeSiKtXitze6UaB9ljI1rwD40iCrdUy/iVp2Btdt
/HkI0E8dLShms84u9vSxgzOWWskXKbhrUjI7+2xhC7hinAwYCIoRO507ozHHgpjx+Vh8GsOPIsW5
b7T187DaELCJzoKvKA0X1z6/V27ydwznpsf/KsKU4zGZWzAjIbko1XV4xUc+ZbdHaL2wH2JIZaRM
jqWNHBJ5fLIWsV21oCIHH769Cgvi7X2s3PedW2OnAbCqSbpqxhdmtTG0rIJWKx/Titxuekg7rJZ0
+vgKOkE67LWuUtF14aHil9gZM5OGuj8RqRNtJa/awMn/VeUUfl8lKbms3tNImp773SaiYMDldZ/8
dOlGPk82n1t0XRaKoKC/ov7JhdgryUNLSh6Rx7BQs7VDlsGWBDY3RoLwenIwycsOC20YxTTPYElE
A0AnoyD56fRWtah7BWjqcOWGCxlDc4XUdY84L1vps6JqpDxn+SSMqr4L0cwsE3vMBeQh1CTsOvnx
UPSus1+C7zV4iox3D/tMJCBbuO30hw0EyIlpufMYN6c+8WjcIv0qrIofUEqkCqSksVYWUx6HiKwf
oTbtAvjZdft1QFXGD1uzpDDhfQbEVFHSVWNkBEa5IjMG5gqI85njcKoxSb4st26D8vYy3+RS3WpE
RyJcr9T7AcJlJSv9OPfHrNwGz4KHA/Wvog35+7hZ1IBNoYIAnBWjDmCPhSpLXjveGfOk2ToIJpQp
avcJmS4vIf5i/dWK4rV0di5CuQhPNJSwoM5KzfMoLRHKmjj2eNzW3x3rjJJkY+6qpCqCgB7GHT3f
NBckaGF6bAqc1pzzeR/kSe4iU+smBiEHI2IPP/cGUJmDkLDpZ6MKIXS9jAiVIA51Y+rQbIcKUp6W
m9/JFjYn8+6X9Gcl8mupUgslp9wNpaxOjLphHEaZUe4aV952z7Mq53tALuw7xaUYlBbtr4sPwPmD
9rO+zp55/cCAjMGoVnW5jiqWsB3ofW4dJzVOXkI+ssyM0jZxPJs3FIjYjlQ12ax+a1U6xS789gjB
LBxNd7ofohSoBZuwjOvsrXZIielFEy64268oeR/IB8deWrpXEEH4F5VX0zIVx01diJXVReMd02fu
6D7TXkdUOKgjAtzNSTJv2P3XMKsYcxxP9mS7WKlEvRLafybVdoVbLwtYnyFyBdeBg0U4ZExdCP2S
gFtbP16dE1UwLOr8/Eum3sbJadV0023fqb9ufl62Mb2n62misJBk+AVqBxvWVsRuLoOa6oa4t0yw
O+Sb+8fr2oYZcsgXmYZwMb8yEugbaOIbd9ionCgpc1q8CE5DjGXsBGYnxfgJxqDBi6SjUuivEmUE
KabqQT6+6Nl3/kowGmy+Q6P7T2dp1jSc19Ovl3LH6IiVIw0cDm4A8rIORzkWk/csYhoWM94bM7wy
7TISMNTEfb1QCigkG6WMB1jazECkpxwYzAjUkDeoygBi+O25KGRfOUa2FuihaZa3A9RcKpVK7dUI
RGeRUpGrue8ZkXsjBvMhxQafc2VQNGpZTT6zoTvdSzaghgYSAiGwBKFwIZaM0J+Yx8q0DR0yeyh1
3Jny5e0vn7FVgIewTKJO274MHwqc6aPvj73h+Fslnpt4ozKYbtRBMGdmZD+k3y1YylssOIa3tkRk
bmu0Ml8/TGMqFPQVShI6241mEW5e34XlEZwMp3ysMVX/M8255UBzQTvl//xSh3SKU8ujGCWkrzyc
DNeEONFUBZLzXWzZX9OAB2ooJuirsk8PvKIIWbjBMOxXaBgSfI2D1rSghGfDHUfOAM4wFJM0VcA+
oiJAHhr2bjafu54RJe37cTyDQGzPgD4k8OTQRHAVhbU7Q4mzuOZWzi2FTd0FY3iou8so7udvscSA
xzb+dQdSPV0kVGOiDUw6Ge1MDcnR66cNKZCuM5AZt/Q3rGbWCzsYvLoS+aWMsTB3tKT9A37eYrXx
nUVClwQIQr6syl4vjT4rjpHagIFe5RxjhjJufb0kfd0U/sT21cgAe3rAhbo6lrBn5tFmrfbgmc40
yijVh1ASxC99D09FdkKepzs3EEv9lhwVp8ennxImd//8yxytxehPmFLSo1JuMEZw2oBww6xRSJae
fHi1t1XxhgD21H3ecHxRLyEVLH/hbjbxFb4XeMYi4WvmYxbF3IOKUEPTVfFBDZhwORFHW1QBo6lV
vZruqXBzsXsBP5dJWW5QG40Ngz9s7C3gDeB7+U9xoJ2LMqixi2IKIjb0L2MIRx7Vly7+K3/h6zaC
5o3RV/vJmCC59yUivv1peq0urOlfa6Hm01ki689geD7JuzVGO4itRN/diUov+q4osK0BpUBEwUgY
I+z9D6hSFPoBJd3he8aaeo+OoLRNsR198F4IaHlkCH+b8dOMjo0DjLPYfN4AErBVE5/IMcrj+6kP
SH9zyJYW+aYeFceiBWbXjdKGfMsB4fddgdfQ4N+hx2aDqr7qnaD5u1aHvf7iy0XaHEvTXcA/wzGR
xyhIK+o+Pd3BOndr70cbItzBeVVpK4j4hON6P27U+f3WOhazdNiaP39kLvUD6RxiJuzwJ92uJPYk
ytHYYgDwc4JLFtpn03hKSj7b4F7hWsmLmS81qtNSGNsJQqXv8iVrpoM3DBcOxxL8EMc5jiHqnhUS
naZWDqCKN6C0qSDVc64wcwx/0TZVmzsFuzYaPNxMWy6+HYQ2hl1VQjMSsXCJ98XShP3YMp50ZJzY
G07w2zQUw4JOqWrvJuyQaq9g+hm0NIqq01HK7KjoyCC2rzmORPhhHCq3Eu6vlXdsGcoVda5duDDD
DouHcuRkxsLcEkutTH+r+XGiJGb3DMLe8UDNUHxc3rB6B59Guam4wuenB/feigb9QSQ1E62Xggee
Wiy6To9kNqramdcj5P04DQCcC4i4g7nXFXJjTH8kTANXfRZdklWd7wfLFMzdp2zK17GoWQpxNgcp
hm3r2C77XlNtuf/3XZ3YdHTbfKOXngTuTQzE2PW/2Wcn+RaAj4kM1oa0lvOoaACuss+6OGDNfSwb
wNzh4cOEgC4x8DiNNvjl4qtvHjbQ0TPKSWEW72WJGMZaEysYiPy0sLBwgY3k2+wmPAfkb6pTO5TC
+yhBBStftThy3twf+lLUWaszC4T/flmRTk/0EIe3b7rwunnYxAL5wiYfgSYtvqFgC/MrGoDC9ILn
G7UsVY5MrMUiS7BHuGEOleT0kwyzbB1xkfbgqBUh9McINN5kTV9Dgg1AxIVHpPXVcM6mv++M8uMd
BGsmSLosd3R0QvCL95xO/foskw+AvY2yXYfe6YZ1Ir13KYI6tky6yFVYE3YTRlDjAcRjGmQDlHP6
s7yp7/S9QiZP07QPdgoytAOD0kZS/5GxTw+NOs8ku2XltM9yvXTk88wgkB3gc0E7iNzrskPvp87P
tYniwDPGZIguXTgsiOeQU54iM9A+zqksiu2BTKnOq2YrKTJaoLkv5VtLBbn6ZQ+Sq0Yc0whLHQtM
fuBSthn2c2e3cpZdcGTVXgRYZBApR3we9MSkxqjhG55QzX3V3tP++xGHcz7l2315KKcODQy9XPtQ
pyh4GATS4MXuJtDl0XlAzsMnmVVN7BqLvm/EFSdF9NfWejZSzlV89mE0Ej8oqlI6SqJaGPZRwS5n
oOtQAEzXSXPYdDsiRaOwvlPmrfi9TfwwIxLBQYkPMc7zSp1jQNI2Z53nm9ptbp70pRXzpZazEM++
+sRnJhwlQqWl33pBuSWXT24of5+M0BxGr/mdF3S7rvrXxZt1u7tYBo/P9uiA2PYdRM7Z8JwDtNNY
NLuYYhbqw6eESkOs4ueJ8BKRQMkPj0vNP3KAXJdm4vuN5Yp0HbnvSqJ+dTeABP5eO0zStaLkM4lj
eyiVmpLH/8rHMsa8Fx7Yl8tlNUKS8ZgltIsasQkUDNNcSIn8dvPCBURIrIkxqiXz5uTrDytiahJG
8e3YacElkTd2QFeQuDH2PlvTQ1DCrNhrC40mKx3DbAV0NhHh7Y29b+BpuVI/mszl8eYUrZ2MO/Wx
v63MGL5IdYyDIgUKBPa2UUGadq1EgWssX5/JOa/KDOAsMCHunqPCUEEN4+7JvVnrVp85YdwBigY0
is+6zVjKnoFWfsnfejrf2grCSBjKyhNfSwYb4NVdJOk1COHysO+zagYQtvVaYsxFMHRKYhIIMCI3
Ik4ZxL324FHP/vfh56E1+8Tf8VQlmz6L0IHj6+nuJQaXNMhgxQyqasec3RoBUwqYbqXM9I+9WWqs
yKcMHVztoN+dul1gm0dR6BtGc/C9c9tL/EMdHPnorEgQ0FNqdrZY2bxvpOBh403ryH+4sTfYj85j
D111BtYJ/AZkj4hp2T4ohOTSV8zsTIB336EYZ7x2yM8e9RR71PLk2+izj11LhAr34OdwCRM9JaxX
ylUTd2FhQgTeNPJTDWv+VNfPX9R6xVw6VXQMKuWYcoi02++FeH7JiwJrFmObvwZ0Sox1TcqeMfPD
KyB+2bo53Jh2jxk+fy+UZtIi6UaEO7apicUanrtfBXoAEbvYwkAWbtZEI/OPeiN7AJBMwv+g1MK7
h++8C8m8PilLFn1P7BgBZWjEgP3MVcHGgpH8v5vieQfCO8KpyovWK3+zbxaLaBidNNBRGDSW1un4
nUEC3c31MnxoM5KCGJBl7cnZBxBYJizNgPZfdYDMzAmOG/ZlsAjXSh2Dc2zGx/aEIayTPg0AICPD
l/0dE8koijJq/B68rLqgLeRHe9bgUZGXRLMfqC3KJK3oq/r7lbYSfEvvAQoo3e6R7yPxF53Ybt6y
qOOuEjJPhqD6ZpXFIDUPHkw+9vOiUFIz6GWtg3OFqr0gbvXUcMqaeoQM0lKAk9shX7uxIorZUtcV
w4jXsmbw4wNTsvIwR6mFdUpWSb7t1TH7AjEKDnRCMp/6zf8N0pS1A0q3ngdo8rseY20ViTzDUuRz
GtZDeLmyUxpaf/4OoOooe21xD+BLEjkOAU2C0gYJ3SnYVXbyhZ/nyVdRD8+ph3Xgp850egrODQZE
90Aw+aV6EJ3wYjaMn7otcB64lBd0SdJfbzCDO/g6cxoQ3BWynIL098uViRaysdkzFquAnac8H9f4
fO+1HJ0uByPi1AQLUmEUa+irKFsUDFpo0cwlHuqhEZy2dPGKMqIFfn4nQHZqRu+1lWMuMQTWqlCl
yTr4lvjHmKsIK5Clf2zX2ToekJMWLIJlsdvMzv1L3d69Uc7+RVQi0uMMe9KdbEDGgAVC/6xkDZpR
F5pviVOke5O3xDAwWCiDXWnlD0GyL0mL6raguzU+BNfA4xO1KVO85DtVyn5FxNe7iIf38oeX7ogx
H2fvk765AUww9eJ71v9sOtF0U6OO2MkXQ4t9iaJwrXXcx9NaNNsvqBuH7JfHgNDk6GcsgqKt1c/a
ohUETMJofvk02+hh8eOWPOGFDvoRD0gpYn/CdiuP1IDCKsCH2m8DThu0RZNx7cG21BtpyxDbV2qH
unE1BScaCil1K5p/umWzgoAwhvNOyz6tYxPsXhlX5nRHF0PBgbRogdvTxW/3TKLYqUvE3bpXp8RB
rBmtN0iV6m/w3yA8x8A+1nS3exmTLmCHHQlk6SZaIllcdP1W6mSDZIA1ogCu9RT8ELpNvcM5Yz0v
iF00Pf4Jr9TQvtms8OcgnAmjLlpFU1Y1CsmxYaWRoSvzw1Dr4Bz+FHky1d58gnVkzftiskIGXRAJ
ZlKt4ArA3W7SppOk0HdlPCfMdXVJwkicQPDptGbs5Y3r+F8aiX4v4NeTtDd2+U9PuJpRu4e3Lf0n
uSeIGgjBwl9kbhXf+4hOv0KorVM0F5bmDtTNj4XxjDDob/ZNXGPmererBOONEiXnTA1ZarnHQoNW
6boMzU5bz3rLJe+mRCWBZeNTP9PEjAAOEQDF6q82FslRySKcbij1TWqy8zMloA5vdyDW7kVdXlBt
L9JBSkA9QiIUsWsYMt/j9zj9pv+JZ92wgj7AjQASDG22CyUfJ2iQW4Uq2OUjrzZFm3s+71uC+5xL
IzuYY48Vb7V1hkZAMrrtpG7ydqHFuJVGTEaehJWE87SN48tS466J8uQNUnq0tHUk2tAbGEWzjLhv
Alld8uP9H7Q3aX95b0AdzXP8GZhO4WtdDF4bGDD0o+5l6TshO6akSxpXDwssTszYcRzoEWoXeWhN
Vi8YNOaiACR9jUb4KaW4qPAcSqgd/YXd8WCqaE5AWqrQtddryriPomODS05zvg8Z/QbVkM+/dkM/
YIy2w36FBgGRlAC1wO0R74xBJpoyg9l46c6KAckj6/QsrakXi/R3Zvef6t4Uvls0umtb6t/wuCdH
iemeEg0Q2vc/nMjbbwn7DBO2rehQ0XCOORZ+osdD12A/KiXjHi1L2a4LTHthCgbtUZiGjmSYUxTQ
cWJgqHeOJ57kxj33Cf3wPcb8tswoDvlVjwjaYhgaNvIf+VzvrSPkcGsNHP71o8pPjN+TMsLhKkMl
OEZFcy4D05zNoBQ/K/0lwkSMrOR6MknlX/5sfxKWeSqgA6W1+hzTZverA0eEoF3TQtVzJubLwH6s
YXF8cI0BakV3BLLfyT0SxspLUXs9uG5F/g4wZy0u3NXYhd/e3X3gnfl9bRcqJYSMy0D5SZKQh44O
MZhcOdfbgwy7xdp464Xbm+gCdQaV3zHkNbMcI4DNQ27aHaACLDCORsefOKJEdhXLiqHUtsV9A18E
UbWfQagpbGRkiny2F4FY5RX1rtlN9rMb6AKZieAwGEoRYKSkX2l1dPnwyvSvuKEWjhLsqJuJuHFJ
F5NudhR6ie6mDAfLl63XbAQgd1S2kUWoxuzwxTjJNNvJ3OPfAidcPzISzmM9kOl5k0RYL+AGtayE
797Pw4Qh+pawnQJFzkhS12ZWAfh8Kg/0mWOgP3GhkdOJl6oU0+etd1qoAB6Lgk5uS5OIGm4vBR+7
+dJKwDs0kKzGU/hwSceoUPrykW8CfEC9SJe9LHGiEWLUeItnqPxZSzCMJ6ohD0Io/4mIZepr4Q2k
sHq5mkOQK3Fz6+yc7YR4vOBQmbiRj+biBgN7z0K5IZyXjU400nyK7LhQz/fBCvJ4+V4pEWeuG1pV
PnXZ4ZrZ/E1crNJDYQT+/MfxROZHKk3HhsOwMWg27FqQMCrci0VGswa6kEbuwoVm3ycNJioF1Dcc
rCjXtmsrQUuyECMocYLxP0Z4PoVnS7hjpypOfEeXYsKhdjzHF1s0unWg19GBBaz2grpAFcNeTrWw
nIyahs3tpRHbv2HCIVXLvMXwjcV2ARR9Olkpy2amr2ugYBY8y/4JqvH6PU1JfuthijnMIouGkRAh
HbTNNBtA1VG82Z79AwD1+UiydpPWV1QaG5bKv/IGVYbbZa3UQLrrwuJmYM/9iFlZwixFE/qz3h4Z
PW0mYIynTjpfxNYQoBSwK2L3DDAi48G961tdn6M7smTaje7xA0gDie9dnx/Fze6W+CHiCtYPB2pK
eFHtty5pAjoYBr5KwfBxVAriVFJU+IO5Ey3E4iQLQLv3PUzv9OFQt7BRuNE6zsyOCW7akLe0g6Tf
nK88mvxtjOmDMnPQ3u5jFbayl83lhc2QSOgMMaNMUs1eVBCrL2AXMK4sM06M9r/g91ADuoqCadRy
kADNICFm4Zc3CO66ctXxpSYwZT+WA7UTb2sxLbZ7dSdkGliTIhXGsAbbdByf5Fx9vCIDSRTxo/0F
Rct+MqBx9PaFS/aC5XeDIyUAWBgHLm/fTYEBpWeCgcElP1C5MMinaiI6zamx8dUMWFCa0HxhKH3S
BnB3nZHlQFU2pcyULWMmC5gX8w6jcKpMFg1hEIhAvKozBSaP1oDvLBYkayv5M4FGtsrYugP16OzR
oXDqDszpEjn8ut+vnvj/QJ35QmpfcMySef6vqQTs8JA8I0dMCG2gvWHDpk5K4XY7fFwkjC/6mlZG
uJp0yxhiWssKhoyyhH1b/cPbE4cBymgPfyUeN/TRJ0Rov2DksIIC4iS9qq5i6IWeamzwuDM0v+kn
d9mRHOKXgu7v14Ross03zkwlN+XkxY2b0ptnrSDLCkmkyDQocMKwmlWwi68Mmu2J703qpv9/T+4l
izV4SdLi88PgfZceaQ195CrL4+fsCKjAvRSiD3LQeo28VfprT7YQgPcKlXf8wN7d2lXz9cZoJ5iP
el9EPe1N6khV73lolDWYEnQBRu68rDqfW095tf6KQbTUjeD2Dp59f3u3I+Yj81JlQcdMb0qSFlMj
UQ4laKsRptj6ZJepVLGtblBmm7YqpAXjeg63pOS8yllMj6yXZAJu7K8p5dwi0QfZ1pJbQKZecA8M
ujhjJRTULAC//d+gzErdHhFZTiQwCQJGBlaVBJnz27qJkG1yF0F+JLwWwHXrOANwdg9EgVh8Uy7b
2CVRtUFX+QtPwhzbzxxLBORWN9yzlRMlvXYLlw1f0cGhsG4avuHNtU5OlaDSiL4K7uuGhg7VeEhP
fyLCnqwIqhWieB3ciTigIyf0r+yphimWfaTvWS++kRLGllP/Qa4tst8jhqnLxvTBrHNSuDI27PFv
MaoxweVs4HXL6ohZl8A0/wF1edd2woaAk0au7BNvoiAGtAmGNr2OkRSq6SbDj56F8YO/AksJ+7ux
nUPOXKnwjtJr9zSxZgi838xiJL2sBKHYiO0fEOmRIs3uli1Udjyalpmb/ZvxjM4f1uOqZdk16ap2
GySdf0AismT/QlMhYp1fjLTq4kRV6gy7UFlRVq1N5H0daaoJ2OjwzEBHhgiDYj1uJCkmlQN9mkLG
I8qXSm8KKOzCnqVvt0fuzC9JtUVRE38PSs7ZG5VU5Fbbn/OOVS2yk4WrEBNoUAfQ0FyRyWa+AqNG
TTfWx8BhXVxXITQSlZ9O+CcMpw33l6zIBH5LvaHryFsO450+mT1iez7AJkqTRCPQHXz9EJbnDA51
NbrEoEeBpCdNaZha2YE0lszprY2AbQiq/5kR+WxGLcVGEfmHAZiCIx7Fx+aIo2y1gEOW1DUtkrZI
X1RygwGU6fvJ1SvJ2LlsCBaT1lX2rCWud2G9P/2ke6JNj4asmvTQaswt6atsKgFMBAP0+o/KsqMi
GYtN4+c10jQTbLlg1XDty1hrvb1uv30mLT81HcWvhnnlr6cV74HXI+ij//Bifs1PuUV7tgGQDKJe
S1rIFcE04NMJQJlxCCmPydn88lx96zYXs1/gHLG30BNFykfF3jEMyQeVgOuJQpASpSs6Upr9Cfm0
QifnBXlxBh1M62mVdb+23eHNkzG7ppzBCc4ZTx97ap9YWgGHdGvepePyQOB4DO9xKzDu3YLt/lAY
Mj0K7Xfdo9FYjn52dCBMMvayO/RFf5p3AjHyqXojNy3wlXIdRzk/rKC2s53Dj+OH0oVH6J5z0n81
CoiSuB2kPeVh201J+29L6r6O5E7jgGoqNn9/3Qjsv8UpM9lqp71E4vdD7U/NIgVglgjdlTihnjzZ
KjG3iEqRZIFvUpIrkgfKYvqYhgHI8klOv9TKfknp8U3jBhcG2OSO/TW6emSC4B0jHQGzWYBvQTan
49tWiZ2jKAGJulckCN7hAJ8PlDFTWTERBjC3gwnfLkJghj1MZttSrNVDkmjNIxw3m41Vg674PA+5
49keWIM1SL2Gjs581bPZYTMOrzwwqJ9J5ef1mPHumUQnsBE95b3tyvTi1vcGAyLzYzk7xkLqQS0V
zmWNZpZ+rApscAdLRvWjkoJlCtCwLRCJ0tKIbiF0QGaMiFUXE7sQVADKQL1rHWGVDquhRSq5R8l2
5yFq+sLT5yvFoZrmXncI59lAczX6mn31s/zFUKc9jIQcRhfZKPG4yLAeCxwlVhnczywUeWlnVS7q
FyuobyduT2fxxj4fC4Er5H0pvFDSVmEL5+D87paEydRNj5gwj7mNcqCb4boxkgD4lvpEyUP0TCIk
C2wWNkf2eOer07uZkjozwaxdaYfkjG/9voEhxGmFZt+E5p2AMptcRRMkWNbvXph7/GudYxyBC0zG
Ae5t4M9hUzaVytoYbszSuXzukqa1gprqYKfUE2gnhKUDFUIuAzd2eOl5Kz05U2YG0v42hjnSy/T2
TpufTbVrcpKYTzclJv731F7EF+qFZk26IPMjARDDiwjHGkDsI5wcmY4Ogv78uTZ25TjsRvHJcant
3jMpR6FDC6uut/donAUdYYS0/Dn30UVZC7w073HtqBud2XCrZZD1fVcTujmweQWwWZ4tN9YuH2UU
+hcKw1HNzozM2hDjlhsrcQ8pbJUFVzEx0cQpvxhW/IKFNUe1+9K6fuqdubPOiFaDJNq1wqO5C8P9
fyoUTmzKYpRPKQMMHmJUftE22+ITjVo5wRy3hNnFbpB8fQLGStxGCWzAK40O8I7i407Wh+EiG9uL
GKyXa23ZiUdZESQniNNjQiW+UsdHZIBEFlmk20IeVWO7FJJQF0DXA23p28aHqlu90eITeYN/q+5w
jsPRwgOlsZLrx4Pgp+PdEbOewrN7EYP9PdqowU8SYwmsxGZtMz6L3wZPYjchjRsy/RIZiAy370Rr
uKtxB0FMx/blCeBEE8x6UPk7rMGJrq90J2MT3JxN9EMMAkTaAl7DmB2e2J9vKh1WFP3S/btp84Jx
Dg3vz0ALUq/JSNrmfTYLFYO5Ijek/O9wU0eWDz6HFOtyDDpfV5Hl8YfoqHU/aW0st6PkhD8WX/3G
sMJYUqp225imaqWWJdwp3alVFl8T4/LlL9wRG088jvdH+ByDJ3u6EnVdDBKN/p7Cy8KHa7Gl/TaX
O3PHYBDOvcCxkJZ8EBEHaEsm8ByNrT0gM2tTU5Wg9h0kfxyIfWEww2xSAli054fEiF1qf+y13Gj0
3PEriNKh3W05zmn8hJmQ4/ixTPLBjSL5ByfsAdVUBaCZmIpLFhkaMgiOIz6l9pBkfy5GJyV0PyC6
vDMud6atR8/moL4v+vhhXbXNSWNXK8bivVKXe7q9L/TAJngTCYIZASlLjXoNptLR9vuGxnxcz8xD
rvPM5l2gSRGFT2iCT8QjtcFbms1JTWc/sOC9ZIyXDcxhv8sUOQHzc6SCc3dETegQm3VdqZ7SOa4o
5y+w7VIC4hsPMOawN+4P0JOJTLTP3vAwoaxzspSfefhieNs4JTj+ZwGKuYKnHODgb/2R6uiGPL0P
Ll7Kz25+TOT6wOHwlBFYXmisdQciu3Y/cMB66MeHU5lmEm6JYf/4BlnkiU1LlhJJEHtSspvsZbSi
jvXxNPqV+CiwXM32uDlMfFZm3AlOCjBsP7HzF+EFebCoU7zG+99kgFeBTXqAGrIKbHqV+E8t+uR8
CRvlTpIcPBSSymbl0I+tUIbftXeOwigM74KFvXMi+nrCAdMXSGWjDR8qNdRSdeiuIImJkNhcyxrt
KWVwc0BIB3/4/zvCxkfnBApboDkQH89onZflHFiGXVH46+X7EtnxTRXvyOpA87gGSOtyaP7QfPZ1
w1CQQCnyeDeGh9CppsRqdMKsrrpq4AbCB0X0zdinQ8aVoJw2jKBaolrOUEruF6kDpcWI2K2Ek8I+
AT93u/LadkjW7fED97BsXDRWI/nZoSqpPe3RVn+ytbb5BI3J9CdwvOaEewiK7IrGyAVadjg/BXG0
9uqc2kaJSptkhaO7HArufw+3K5t7e5h8GyUEPHyFz+YplBViyNilH9e/I7tp3b+zV9T6AzK1cTxm
A7ZjJxDlt6ZK0eGRlGYoXeHf1PVaHIU/K8eQdh/Boe3oEjK2/0Rc7CvlzEvRyf2fopAdIhd1Cmm6
M9DJb4pAuffqS9J0/eCrCJt2Q4rhR3J0O13gxJzVEcCF08TkibHpSUxnKdhqwPrYlxlsL0IvcXi6
XyWSJ3n0IRDazPGga8hD8WCsLqHOmr9ngJa36l0qmFhtexs8g8DUZtWABEOsc8PKtryVuC2TSgK0
JRLuDfUeC4phipX6E6OKPMIGyB5zADTxsZClAM5Je+5klMV1PqqAE070alrYkCHpn2GUuB02H44m
gsTKJ7Dkd42LIW/R4YK7RJszI0/W6Id0vytrsdmF4H9XFQn2bo2sJyTQygTjO2Cb9ESTTOWPGPwK
BAevxqdAhxjzFDulswh3AJlgPqjhfQmwt+TSa8BuRbbFH0JLsXEHSDjXw4K/bwwI7GBOM/rOEpyk
NfRHvA9m8RjJBAKFvctD4Ne5w/+sd37bgFJgAB5mhsCNtNZT53XtMkoKw4om1Dws0oczXupqYy+R
r3lOi1+8N+K8GLOcV5SgSHqwRQscMH6UEwswvt3FxpdHGb5ejLXoAGMiFLPUVL1RZ5FpkaZnrSs+
QaEPElBasTRWo2XntWTEIconFLGKHolz2UdqDhDpXyQbt0GWISEkDXzovsyrFRGWu8+SL/oaDL5l
04HjMnhZoOMT8J2tQIieR+5qXxQiuv6P/lL+78cMtPKRwoEKbWdV+ZNUbQGvCtGJFARl+sIJ1siZ
KcgSAItH+1hffo1ypiKZf+rvLnQIQaN/kNys+oFXywKtQhFUz8qFjsO+VGZpgC1RbsO3/gJ7vTqX
SgpXYfkDCGz9qxJdt7ROjRNUX0rH6NPwYuketsVkrq43q+jTlF7hvyaZpV9r+ZL+IzX3elHp68uj
ywuYF9mlTcZtgft2Y8tJy/5ljoqLkCVWY8t2eLLK4XgMDKsSiABRQYzrd8QLPxahaX3ZZT9/SBuT
CGcjMRUBYjZHqSOkxClOUYOEvzJNVGAVHpRvFM8a7y3pmvhYChHbQxXviUi/mR8wjJp1woGLCpc1
QQWqRtjM/ZcSB8rzmq6b99O3rzeIs0Un6GT+U5khQz238norsFHRvGwK8hFDTf0VWDy/HD3A4PSL
5lfvFZ2ukBRJ3oDhxZ9Cq6uwisEB05UeoWjkWuYctTLTE9THYcUGxN5XqeQ5Mo45E/YI9Wti4CKX
usoXHZlZoSp+qp6MfwU7ZDFhrK3I1OPaieDSmufN9oSE9ZUtY7auDK+mOFjFrqwne2WvJ5Luv1zx
dsF7DAKYI3t7+/FxRB43u/OHKZrHob74zlYsrU8bWiiUm1LqCqWfV6opLyPGFCZaTDZCJTtT2v6i
FbxEFZAInh2XOV7sre8DuiL2g/N8Oet2Fht2/VCYe6v+q4z8ON3771KcT1VuTtxjka8HB0IFTAtx
YHgkx/OBEDe8FNArZutDtxK2uVA9dAzHM31PPHvqMktXsgKUWkx1+Ps0kF3Ql55KN2c0al7/9+sw
m4PBp6wSywroTXzr2YWby/lzTlnZKUzlLw3QxO60u1PlU3Ra4eYC1nVultdvMByI/lr2oEQOHg4d
PB45eDkUCFy+LtQE6FKVMedBUhXwyThqMGLEVYVnc3Bi4O/vCpt+hLPtuSYYmk5RUccym7iaOhoV
FHwZSTAsOFn1Fu2T2KhmnNRmGwfwmTcBqBVVXMgjRZ0H4GxuxoqmSahBVZHE9MlYMlTROYtLgvUi
S5OBNXh7Aq/c7WzVoQufY0ZMq/hEACI9jgaO/9tan/z6VrlUAGKmvwz0E2QRDV+iotHWT6QzEoU/
Gwx+3SN1RqSzj0WNTsbcL+f8Wy8jVRSMkfAplnKOESkeoK1ble8OJHxDTrPRYFH9v2BLC8bjOUTO
kmvWmL7P1xKe3Qh2dEitbr48QjiyCTpkIHSQRNfw0gA7hqMBx4Dbzi8hBgcueQy3IV4W3hRgkZ88
RN4BL6NHijDowreEnS99eO2d74YG9JkqyRmu/IpDRo0IKXuER/aixx3lW3i40qX7IubkgHwJUexE
l8RuU6gqXIHCtH/q0gIpGKd/Mz/28y0t4b4Kq+sGvKF6LOb5H9bKwTYJpWgwR3BKkLnHPyxENgk6
M0yJfdmZ/+0KNEOABHO3qf42aE+84Cr+rqrAAL8icLCTPkgpk5FA8XOxuIyyrItA93a6PG9/JVdR
AzxyHEYG090LGW45/Tg5353Haqv0usp8sWa/OmfsYkS7IF9TyjD+NbhYl0DBUqtpfiqJyP//iNnm
zr4Pwl338aoR3+rhkWj3UfyVMtieqa/G5RXQGiVfOjfJUvMZRxMPZ1D686lSM/UfMHbpMocC4T6l
NRLoP+QQKYnnEIaHaroKGdeZwWksAxHEUAIHCOm4dxqyj/8BG38eUTuGBwWJ7/XnUdQwcldMw6D6
NWzRFeOHULiJMrkn0zBpn8Rd2ixeRsdVc+YaJ2RWPsQkN/dCX7FKfswQrKVoTKN5d7Dj6i8aLikR
+i9P6OShNfBQTwcmIgnuzIpzVAiyDSA/9HeMT1gTvl1uGdeA/2NAzKSxYVlSzzRU76Tl5+hsDySO
gyVz5c4SNfOm4XIQwU7i5CTsBI/3U2RvHrPx0KqjE6UC5ZNadfxNML+4z45BSGSRm6uJgIKT8PzP
J9qZRsWEgYpLdKLUgPuDsWaJtKeL+qcAMn0Crv2Tn7M7f4UilD9geuiIBB93FgDTXe71GGsMOr1N
Na+a+IibEbZLc6NedSpMIzZabPS0qlhyWlC9qv7WW0eou0Ecom5RjArxdyGPuG02jmHhEGg+rSsU
rNvxtaq+4zoMQl9LZmfLv+szazAzrKbXhbjdbDeb6VgryUdu9gTH2WjVbZk57w6+qJgoqeNyPqFP
pgHhl8zMurN3T4svT1n/aZs9CrQ3upRlj9Thid6xJYmWfDZWO2houvtYgK5jl3oo+gv3JaL+q1LW
U1gzv/OAiCoepqi8SUz+2RZg3aUb1fZwj2PsxRmd8O9ovHRUmDL0KWW9cw0k29GyklwQDy5ubLQX
ANTQm7bf8OcI26cZP36m8pQFVn7J+2gsi6ExV6t+tPSqJsqsF27gQTjUrP0MISiixJ25cGgQF0V3
ZvW6ftc/WvhDrXCpbVlRA9gyd4bsGrNhLaU3/oaVDp4zEiHj3hloMuyTiXl0GTHs0Fbd6mwAaiLj
BNW9QqBnzg96DM9z0b6Q3eT1tdIskBvGvNYrjKECQqH4TCzf3dNaFIxg/kDftPP6WH7dTmq30sQK
WNV9QDJmIE2Mc0ekyyj/GA7PoMhqx+kCz60zOhXTQ1KV7azt3Yx6Vkt/hqiKCWcAx88lZlZfbxlI
sK64WyJqcPWr0XSCtKz2hZ8Rgr+JkzrzXgmzPVXGpaasFND27hCdu3FLJrAJtvEIjAuZiuqUPRN5
ZcQB1AZPl7F7b3tCb9MLidathUkzWFLOrpAN153/otd1/7ONkfxVoWS3X1iKGB5HSMPmsb2GvaOJ
BoOvC8zb0rwGDkth3gjoN/5+17P/YAOOjG7Tp8Fh4Y698jquIH+d4DhYT4C856Qv7Al/zVcS7NYh
jjdqQVdOf93Y4ILKVG2OEsUlZEiiLDANX5xfGCQky/pqFg0BsfwPNl/KhlVOFMXhUmnMlilWOabl
nXyDMXNBDWKHv9TjiepceoJ4w5BurkiOJCyyqmflUfa/+9IaPAJnvp/xdnan3N11jZ/oopJRDzKd
FdEHbubI3whNqCnbtOpsscVAAPRmwTImUPytmXwpaoYzfeL6ugm9tHsc2SGy2062n4tDDxZm4WS8
kzfI1yfat/uPF60cb9XcL/X/PnxNm/LTGjWx0hrO8tfgICk1lTIrFbWuSxm9y8f8fWJVQDuDc9de
7zGhYUDU75MSqDQdU1ydRNV3rCB4J6k/eioBZTkfDCvPKK+fO/d/Cc4wiKn7YO30/G5KaA5TABUA
/RGXK1XdzMYO0W1gg5KMpcHIXCGvt1V+6kQZ66WzgHvpHDnhZGOF3IYDndX4DNpHouNEADYggVXy
42fE0dhjgYrRwa3vmIIY6NgdUmcg+f7gGo6s6Rheay5KPRecosGgjliAX7FDxDT3WMEH+ILgNPXX
Pjq0Vh0pEMEjLoZJScWgqe/CwO+M2JABiiqE9hxaw2H6m2ivL9OybgsKxCyMdVMdfH90dsdkgDt+
zftyzBhiLpyCe00w7jH036YEZfMgslIngWuw1oOQSo2rdNbcTfQhOQE5NFGQGF3KWWkoNA4nYIIG
YGrqoslf1PEklII2UwGLlWO7ccaF+tAHXaB6KT2sNnquGvOH/wDvRMK4acjkurHBEW0N4P4jvcP7
qgfUrqvWt7mxbpNWVoXlLZmtC0oNwM6RVUq7fG+83BYwpwjh2SiA787s/hjL42xlLr1toF5QPwLp
OgpSQLWfnn5ylAYRoWO3/tq+7n9eg29SiekkAElMasSWXTNTqdGYXuIHH5MZssDXd93dQEC435NW
VgSwRnQG74itLGo/OoPwGRHkrUSBDaE4g2O28YoJEnake18bDsI0ALQ77KsSQ5PVNMC6+iphS+3n
WQx99gBJRUySWGEz0hDt+iUM/ZhKSDFiWuemT1WgtOn/0xXoT1qEvxFGc9jIpDN5pKaNa1sDnqQE
LXN0XzVucfbyL/pbEMSSzk+hnoCCdNTmaBe3pYUGM48azjwvlYrHF4YBxx997tjV7SxNH1EnLC2y
NLWsi5Sl5v0i5sgBCIMzQq+nh1R0pSGfYSYYooWjfD5pSrqtiw9cwTQxHSacCej8en/BKKcNGH/t
tF/QRlGb3BzF9GJleIqhceSq6d6HvIlMGwbnBuTye0daWG6tW827qIFIg3Rj/K4Y+sGuSlCCGSVO
Rfi8ibPiNX9GvZEOUeGbBZ4OK5tRwP4SBtZI3sVFMVKjGMO15zbE9hgjzb43pdPrhSFUwy8/HXuX
mqPQJy2wtAmZpZAia6asOOZJIfxOCrHSrYZJOniAtiz/kYXHtqJ2V4XuloL/7fGHYj2nqBCsxXFD
tuTtJG53IOXTealbs+naUjz4kDbGxbZ16EUBYeilaLQ6PgVrfLOUIG1eG3kONZ5STwY8qAXj8cA2
qqJY7e213gEw3ebGTjqGLZh94X9XJn8OvR4sR2O2Ucyoi2iK1HI6xOgdbUVEZ08Fok1LJZXLdBW6
ob5S2gThFDD1EIlx8fHA/zkxLhGF1REDg3xxzj+JBPkxG7uHfQuEb0BWYYsyY7hICJfGUEP1N66d
4FvCWBX+txABxOY+SmyXP+Ke5Ec64zXf+h2df6BxI0SPsstefDxrUobQ3AduAXrTnze9QFworp4b
H/b+u5lYFN6v5AwrQp9TTHkW1fetiP92kWM0in+QaexWKLHsN1v2COds/8RNLp73rdlyhrQHtQUU
s2lAm2FdNPjpn8Q4UD09WBKXgysEyFjvxys4qvBAFLCbNp+NiZiDJ2ksEOzBwCuaFkPvNDN564Zg
E0SD6Gj0nM7wX3iwaTgnTHJTHrQJflJbRCbJfFXwZKm5k83gvhPCImto/+FFdjBTlNGflnjBNep1
rmoAjOMH3Y1exmslGLfByDo9AYVkPSlYjCOffyUYaUO0ICP4sjg0yZisB2E1XFYpQhZOyHkm3PCG
shkZbnY1Z6fE/19k/H+0WLQHVD0eiDrdown1AzIK6/EDLHMAVz6U7O6Z4EJXgZk/TfVQOtQ3iNvP
II6iMGrcajsr67fwecJfnVsxSsJVhJsG5kPBOK0rmrEiB8SSuuCaLIXPbczIobth/RN2X7OzxSYH
rG6nh7wtMSuxcoV3bcKydcKgIIkUkBMwkY0Hu1MzRI1Iovkq0WJoahEjP5u7/BTdwV0iO+oQb5Eh
sfA64US2N6PlLOPh+XwRqo5Js0FcC9vMaOimLyoVdBUGtAQ+zNQa7FvLSfwzgNOUsQWpUyHHpMt5
P81Zf0yGJMOApFWP9uZziN3TpUpzWd+/rv3R51AC9xmhP1mn+Xuur7v/ddz2799/LkgXD0w3Cgyj
uOLCk9PXTYnv5V970A7cbtKCwS3avLCghjkmQwqSchhvHOqVB15OcZMnfqYO4z0mk/goDJ5QCwYV
wstktC2LbSlyPkvEROVc+Gy/JzamaAHDTGRVoHB1Sh9DorOmrqtqIiC69YkmMZe7goXvknbX9aym
dvw5rc3I+wUVTsN6ZLq/ZLUrLYA6lc5XTpKDSZfp2Rq2SLAZngt+Dc4XSMoLslmuyWd/kmYf/qlS
nv7T1vOVdy2b0LhgzG+L9ImKEKp5ljk2O9UDiSB24V8xRahLFTOL69b7BCS/hhAXky85IQZp4pSP
X1aCF+gxLfu+sGWmhCf5UXcsOSlRpgEcKFjSvQGh9xMdZyJ1u4ClC5GqlnGyfVAE2RljK5n7qpYP
U+fvxxqBhy8KBGjaJv0/1754MB/cmoj5DneojPoJ4DPTPVjIl7EmP4zolFoc4BvrXjT3C0jOSNIg
/TTwihRPQrh9qlqqZUzI76kJHLp3kGahvRlAXRTK/mNNqJH53JfDjCeG1TJAv6SUxQBBBIPRWLpN
I6P4yCOGm4G58pXM8zOTf4bovmhzsTSIJKQMQdTwc+jKZfwsLxoAFB4L98Hhg+6CMuLRdGg0WXjh
YKGa5rrKe/j08eHUrCl0e5/QFmqZBx5iA8u4f6uRUoPEUbDqH9aXNiGcJLeaNuLLdAFgnz/ZQZ+M
7YQlXiw8xaBGNipuPklP9WrKMY01wT/UN4lf6R314j+4A86Y4TJjirSRHd8TdQ1+t2z8uNcE+TVU
VN+L5v3es3QCSwLY+fS6B0rKxiVsmVvwbdrdcuf7d07fndz9W385w5v4ytkI5uKPPUjxMa65ciru
A4h+mB6JMctBmS3ln/VHG4uZ649MENcysNLB3kXY84jJuwXnCQu/u8PrppV3et5+NbKLw5b04tZ2
s86NdKTcVR07b1hc/hbml7pSpBDThFSCf+Gg2Ob4bRo3MHZNaugfblYnXgIxsGzw/bj0nZP61M46
1rRhS83fsNZSKzwh3St16ujeZuHhGVg75uooekKj9h64mRshSQnNk/HoPWKLPVab4UtYZK1bgo4a
YhSg5/c/q+ArwBMLUzcyKJjleQoWu327R0fcCOCWPr516kBKitpLCX6dKBJ6MJQSmf2hKpv7df0M
bPt31mIFhJo9H2KKnLHr9wMYrSjGmi6wedbFjmTAwX0VMENLpcEKS7B85+uC2zJA0+k+5Kr0/7S8
/g5CiiTtxczGnshmd1qcio3ruqIp4lT0g3Bb7P19KnmseCzhfDDWioElUrc+Tulb2RkqtDoEK0Wl
51LdronCOjctj4l0oZ8cd6pa8ZLDUwExEkw9l3abGe2ppKWl7SLwkdKtTtzcMt3XBx/Yv2eoINep
DjDpFAldondUes+DfOHlxw3M5+20tiw2b2eGo/1UTzvDFR62BiYveWx4Y/xmrCKR49TrPqN01voc
tDCzwowP6W08zyKLhCk0ovXW00uSCdHQwXnDyiq4C1aR0XXTEckKXGeypXtE++7EQAz903UNrKNk
k9ueQ00izYOpE9QwesnNtfhOHh22hwSavgcQS5fbFDPhEYvzueTb8K8yrhgYxTJEpwNbBfE6Q0iO
tyF/SoPE9e8YRJjdEXqI5LzFi9Fp7xuYpzs81+Yezs2DfNq/0E8FWebfDsB5DSttAvkKv2SFrJjc
m/rCFdjzBq5cgkJDd5fO8rEO493FRBrOGR4uipr2M+f5Tspf+DJNcmd6+SU6A7mkYfV/Hrkp33gK
9Vje8gJ5Z16F2gKcjBeBL+wxilvgeZtEwChLm3YXeznHpfleFr8J8R545LfqEPdXKM/1c7V6dTSa
weOSE+51VukZbS6zAglVm+rr5I3nAdlcAkGe84wAdxn9d8ysiorWacVvTqMANPOKUxXjAAi4XcFP
Y/thw5GZ07zxQvtiCVbRxtvDNE31sLYYSOE2XXDeJKp20BYqLNkDu4BVNP/+W5td07tGPcFAPnnm
CF+n9BBslc8V8j5BCKnfvGd9YMyRNQiGd2hOuV6KnfbvaraOOQkOWTEta0f6dKlHG3j6Vj4O3NVa
i6L1svNhQvyCRMIYl3lGpWcAbzlLVvWnErzqPzCYBaLpwWzC2F3WsgepXwlnyB6qI0fzeG3KLphu
AxmfJ2WRNwRZ1arhvC/b5T/zCrYI6ht6t9Z+6tF/LRxuG35/K/U+VeI5nJIk5IeeUqr1fqgmPTBd
I7t88UvGAUh/mRNwPVSWl+wfBMYOmwIN0GPj/7QFsvzJ/sL2020nJMNyGuU0dt/U/ZaF0MTgjA/T
vDKt7kHkgqnIx7/f7cKn9Gn7YBMLRX6Rz0cCb91UDgvFtddbedk+BMkPivnXZyTzYlhDep6SPL02
wBJC4bJMyhFe8tTkYci/Edh+vajc97WrMrGMiI11duLJ8cEhUF1lLOkfASkCJ/CaRv8rbElQDVIc
WScRW6ufJUZAV023B9EEcV/LyDQn5U4SVrvhD0glwpKpNFqd4sqVLbEQP8fU/EPSeLJN+6/QIxEy
UBEFR33k18iVYQaHbof5urnkGxa2rRm7+E+Bl6XELk1IkcjcK2e39vihVkbVxdiO1BdupxUPgu/l
vxDP9FZaCYkkyejhSPEiwFZB6++6DUaMgMdBWtXVtdMCM/3j8vKGLfbzaesvwjK8AARY/EOfeWA4
mEqdhhJr78wpCgkvUu8yB4P9XNLZTmBV4WeuviCo+kwoakel9D1QRMJODtsxbga0VVVuBaDKRJru
U6gs7SN3oqWf5Z1RsCVpWfUKUAvb0DtYfdW4rcPFXkt4J1VAiCJCb3eFQu2lF8ej1BOwA6j6CLqj
OiyCZPK6bYryiGgAFd6k94KtjLyc665aDKycG4tgWLd84hzZ+6m/rOkWOV9MeuuK0vmzodSa8Cb4
nIIXPbu8LU8daYXH4o3kHdb8ywuRkTx3aBBY13u8XxHwsLcwT8u2E5Iqqcu+rg/RElp6HdH05Vj1
sXY0xwVxZVSFaift+rRYXrJYKiXDyAR7pyKXOfmwccoz4lEoyTFxZ2GCDtAbjZGO7J8hYwTetxnv
ZGKu8KYi93t56emLGgb/+mP/uglyaeKwwRSMTl1KVNa2kmFUA6dSpAjsRlPba7eR1mIXud92hOLZ
Lbf7o6w8ljt38tp98/dFYG0DZ+OLGPRCUbnPqo4OvYnQxJK4F5yCdh/kpsMRjYONpNv89fJiUchj
L+2shZNwGzbZwt/7FUe2JMojQzdqY1J7qv5C+qgvJzb+8+dT0h5EIS5r1Ql4y8ZLqAv+SHzI1eVl
6rCSxWTXNka+1qbhVN2b8W98Ifo0ACO+hhaxXdKoNh0zm9sw+Y2XDShNuy5majxGj3yqxX0Da02I
MdAttpZ4AP+Cqr21al9E22gOJ25tYo2VgPpvt0SGAeCx2bX0bkzAzi44IP4DL+UNfgb00Fm3W7wB
0MN/UPInYAgkC9qHAZRooQLEKS/EMN1ZUUJen5TFho4HKGclW7zxjFo0Br8KnC8CQtK1cWaCZZSa
yRUyaFlwzjQgKqiAoNLyHAeYHOcpR8rolE7WDOU90mDBpZJ2VEw3Jj43H3Ai3oQgdQMv30YZm0zH
yIo3oh/iKUiSS4gYwY4beauBSxdHefrJlCuiUx4hkT65NbJoxkPLGIeIXwDHdkNTQUHOtXBQdHR/
GuFHDXXpOQu1NyWpfar/sl0ZQkrVpWJLFbpaX36UQUemUMpafj705Jo5GHZ4Ahnqqy5Y01KmLFv5
h/pNrjfrgeMLAOOs8yvO6HfZOsii+FVX8W09NxKjkSceWOD/j+PoLfOHWvyVD0mG7Rrrra+pLUyL
SFD9cHwhaxyqLQPWL+0zMDnaoHQWR1fTDqVJKWfB166f6QrGeCoonsoxBKI96O3WZZM7LEXFthz2
n72SWaGwwPEUuQNGCl2v55PuukdfHNLmuY9KfHaVlrJYbjXtw9Yxln/oWareFiDPPQUjK7qHQoyj
oOtAOAP8XiyH4qAFlASaUhxdsMbPEM6090cEUIF4N9apUcrLxJea2QyG5VANTX7rdTJnJs2DrdY4
czcSSENQuS9PVNYo5cas2STWnNBART12vVleg5pAJgt5IFGZDqYEJdJmOZBEYlxaUc+5DJlKth5B
4Ufkk7OnY3N+++XabpE4CRCwe3Bq6QlFi9CMopHbUt3qok4vBjaQuHP6Xu2OtsqJJOTAG/uGXWPw
C6cgZCyazjEj1SjTHCJe7IBaZuXoeL1Q8Tnprwl/06A5nF2RpUVsPKYC9uBJDuB0VOu+mL6Dzvba
r4BhoaaVb689Nkmst/nKhlnrO5PasFlFQbmLUNU4fpZXu/ioUmCgiCzDLN1LclQTY4pf4pS2A6+C
AdQEgAAJUxR/yYjSgmCdSKWUAR//yafcu8Bs9N6pwzRrxOdwaM8PrzEY4RBUHx0ultptr7+mbhB/
vO76LE/9ROJhKxjxt0HJrKaEKfIfOveRBlzapggag+pJ2u08V8sqSb4yTlaxuY2uPwmQOk5IAHEX
n+TgiQF899KBqVv0sDm3OO7MPWkdvD7t29oaPtxh3fWLSlAeASfZsrrbGCrPypgM5a74dmo85aMy
4GJq+Sj2foKXY3XaBk6NnQGoPT8LpPX9FeLUjKVGWLqXdE+Ctx4G6+NswEhMZB3xamJDg8li3J28
jBuWVmUYMkoniDiDCam5juVIT4ryI6zw/xpdAgA5ijM3BhJBHeialAJq+Tm2Xg7k7OTY8YJ3NdBX
fR6Udb3t3iIJQgs5Qc5TbFKu2/U2aSYxUSKjLlxBZSE10msvYfhy2jIbolvZp8VOg0kb04L2mfTm
WaEBxRS2c7XIy1/MaRoOs/DyOwxcuWllcc9+ET1g2MLiNHwg6reDl4OfFjfz2zVO31SYUZ7ziBlL
2R3CbL1gIAsVUkJXrHNtC+nC3TInQrsaILKAUcTioS70Zs6oSkOJCREwpsgaOiuim5KPRLNxxWGb
lEzoN7b0ic9HCmEfIa/Mw3suLpltQsZyOImP5PwjrL8DRHSlxozg/aC7nal0E8U1d+ZfG6jk039r
An8YJU25g6ZG6VAf2ziGXIZuOmhI1x/3uEQZuBKG36788iWTMBexR4nt5W7o5w7XeqoeDk1lSQjD
vIqgy9GgOKRbwItoIOA9BEHqwXFyXn/f7lp09lhGfcDzvTB6oAw5lzvvKo//sLCmxhQKB/JAr9kP
qoIQmwMXuxMsIeVQVmnaeBP2iJq2wmFYYPXa8QhnydIFN8OzJHeP9n5gl/6O/nm3E2e9oEZ0TGu6
ChlnnYy+BEXLErshQUFxuD/VlfpG/ZqkK5TDg61ALhzUbi3OCcCoD38GpM0fjtdYc4BtF7A1Qv15
W4Z/W6zI6tOok/UOUWubbOLstTsspKXQQOXz71GcgnNr7Xo8Ial4d2umTgkkJ/IPP1LMDyIPIrSX
tmmmtrS2/4CngbTJsgIL8KzEMjXJk4mPH9i/NBhnRX7qshDIzi1s7P5Xsl2aa+YhW39jzuZys0TH
spDsCRUwfHuYfykN75FDB0bxOlISxzH7+90xnc6kSFM20fFErX2342eMuQxu+8Zoj1bQ+HrgZiYl
ZhFDdhuLg0+YPoH3nEHRh0bbidJgEcnBG17q1+WjrZi9UIevvwL0HaFMuWS76eVTqRQPX/nQGa4L
+c3R8PALRDEb7cgslqA8uGK4qAOaTJLq84aIW+4DXBv/WrZ5PxqYRDj/46aq4fkhIe3Yibk9VG6x
SM7A5Txwn/7Y3Wgfd4G4n94Tgorjg/Iu4Nf56YS3j+tfLxq5sZEhx90LyA0kuJcgoDAKcXhvnY6P
1XN7stxfGcRqk3wOEZcOnB2wgD9NJZfkleZakGa+ohH5JcYVYzQLhhfxP5lzpmwpYD/8CgeHJ3A2
H2tNjXHpmo2/AN2s1z33i7E5yStLKoZW//wGZ2gGtYS26sg2+J9OgV3XnioD42ItRhtCCrjcRKQi
xnTzD5eq/ZhbqqbwlKyRRMat9i1bzl8Kq5LT8iyt3l/R+rzmuGWDqTTHDe+lVwVXxaaCvElayRle
pk8chWtnl2JEYcK5LfyvaJf9tNU+cSVXgSqnC5kkv414Sevgopqf0cd4pxYpS/PgrUGZNtBCwrT5
wJYkpfyO32zipg3mDGtupU/Sd7hoF0tXKki+ZG/OUhg00gljaIpkq3LBPrDqHsSJ346i6LOCD2Pd
NPZTRQLkAwlhnNwiQWyl/tnv8UZUwvulsmXUEKfRP02HxJClTaWk11D35Mbvq/n1W04Z8ECFUTxG
z7fdE5Er1QAjl5PyBXDXaF6EfUNejMn60Ii42PTJOOhDxD0y8sdxgTeBnAA5+cJQhFkQxrycnozO
/W9lnFGfR15mkqBNPmRkO8XyAsj40ED9nys8haKFVpRxkavWbdoApEL3CX0jzqkEpJ1icA99+387
LK/Cv5Ac+qE87NS/ur1kdCGXeIyYprngjrFlM0v4Sk+rd69/uGuIzavq6Ym2iN/olpD/k9bLXM9L
G5uzyy7mZ+2DLJ2H+LBOLcsZZ4Tl2c3lTbF4opEEk1ER4WaIHqNtmEnaX2j9zJxviFobRnHArb8M
rz2hruPsAe1IlSlwEhyXCpza6Hmj4yMPucaTdRzm/XxtTU6L8AO+MA/Z9d7ttoHCwgof2qcfGD5R
MEn1Wo0QJKp9nwFuDREBU7aLYx3reltD+N9FEBwaqHpvB2M7GZ2JU97RKP34lnvsI1F+zsgOaFDH
qSclGwKN6TmVSBwE/qGdT71aFhy38n8E5Ac1fbBa0HAfTh4G2/E+Hx3eVsFstHSMZ/uolY/mq6sY
zvCEqwqseucLE/6u+ldRdQDRSMnCdmKy2caLG9d1a5xFpG+4peSdB8uFmZm7hPGWDVbPuXCgjT1B
d6XkaVvY2cgS2Gnh9lxha0rt7G7UUyz9142TXV5ABceBOm+0zbEFE5wCWEkyjtWCbPX+n8Liza5z
CB2QZNlktOrgFJGKgMwSc7U3yKOQMOcMm1GN7gaSKLDYzsuxh1rtycXpyQeJQCvN/cQHye9yNUWA
4cCdGFJsWTCWU9xW/1SOtHcAZydEhBnHBnddBSdJQZPMd78bYAcDePez6YwD6yL4ZvXzhULNv41W
z0Mr7fxIIJw2obOPQ9m+5wtGnkXLPyrryfy7NnMwpxWxa6C/dORdxSfl52Wv1hLmm5gV6tprJSQL
b8YlnYoP/ykM/HFEd/LLV6BkaXHuToEZ9fdTy+jBW7LQHxCOkrTGphs6ITQruF3o36iE6tAn1Eui
ipzw8A0Tieo00g/ctEcs8hHwn+Q32shNrfDC/wSn/yHmaGFUZYtugZAqL7AZaxPF6FFi17Y6sLrN
O8heXei8U230x5w+6U86puVoxKMLsbWCk/ZsQ4IfdsCl8FQQYfhJi7hw0hSEmqv/Qh6Yz0PtvcW/
Q1sBk9lbrEFf8W1GuG33c81g4N2JKgFJAN/VYKmNFkJ1sfhMswZsP5+NeW3rWBK88EwwT2DqcTSR
LCDrNH094V8i+meT3Ysl43DQPmpY+VmnPlzjb34SrPWspQ/ol9WZlveujvU0Jbj1jlgSl/8K9A5/
6rZxm1jP6f7hYqOsLiXyV7j/QUyUW6ximuM3eghBu4zBNZhmXgIIvAzPwr1MoDSeYtBOzbe/C04A
4CDale9Kn20bjXgS74V40h+2gO1XCQpnn/UEghZLemaG/8E7rhweyewWwuPCl4YHkHwbmdbOEfR6
eNTBtuW4IsJv5mz13yTod1Fs/yeJitNZ0zejz4z5qO77Zb1cQH2yLQXqcz0GokDUdO0GMhU/mhT0
9AdFo9PnWPRc9vNuAf30igk5KlIMK2V8qjumyLc9q65bPIM63qKH+XlYnDme3olHt0O0+l9/wRB5
62wy8TiUvzou6XO5VDJ5/Slgys+mRqCnl1CIHKIH3wbpR4EA9g03gkEWTEjoFXbQBaX1jL6QhZEB
NvKWLPlKiU/7o8Gza3Xt09qeLIm0Iy0ADUy4sSltBo3prrXWHaWDHg7CZrJUHS2F5QwZHt+paxll
kjFqaCgcx24ekhJ7KHIpBpx0JxXwnuAyVCHJRC48wpE2ijZX9r8bdPtlkHwNKhEh2jxEE6WizVOT
GYj4G4jq2jIVD8hw24vZsdntk3RX977HpaqU9FBst4hZ+xCS/9BclR41siHAnwxOFsIoQONXTMSa
rwegUyHd9FKYVc2eh6qQiSQstCklLrrSONK3BFCEBfy8z/LHd9LU3KbKSkdo/oPiLpLyNJULTXxN
LRADtY0kE341XvJnC8iF7PDACrCQGvvYMuDGB3V3aRA/9R2xhud8fKrwa/bfzT0T8HZkdG2Fls7r
69CiBXRbbW8xXBInjZV+uNMgj2IlDu974V3rEO4elESE6AuTiV/eX1XCIedvPhQWcWirMhlDcC6M
IzCZH9YhSres7vPILDboWALhbYK9Yr06W9frsedhO8dsOMhh9ol5Icl4HU9DfIrxHRn6vMsD+pYA
OmhI5PCm3Bba0JR1kXshBdjcp7wMm4rJdTCDhLTxQrhVp2DG3xIBK8jHsNq0jSfo8KpBQOxCDo4w
ddV2wJvmh4oys+yiJMsaIplYbKXB8S0M5UNnVofecE2mX0netRmpO2zt2dq4cy1AVJu/+fHFeWAa
LCH4YlMAiR2Ul6axRly65yyDaW75sG4WwHDRJPxcmZ2VZok5TOFR9ARtYajH1udb6EEX0S1POpMk
ZTjZVlD5VBTosPhnndS/nXxhnL7QJwZdTu0xJvVidm7nwPg6VcqlWM8S3Nxl+PNApWXn8OnWDaE4
kch6UneOhCyK37YK26EJcvg+xEsh12HWUC2nyHPh1fdSLzpchMKcV5g13+gtIfpH+rgsvpeNZUZu
0nvEEi6TYXGmdyJLcd5upf7iCDmGabF1GqFSo6ngJBBmqkH916oYnMiYetZ7qmd7RAHXcYGXXMrY
yx6NbWKBdew7pH4RN9EqAM464+ojlxroJbG366w6CbrCoPr2/sMnRQzyfuLyscaGN/b+PHuAL9Ti
yDuMCz9sl2yy29rQrSjE/rFwKH2E6G58v+Fi3Tz7i6TJOzVbKa+HxvSNwKuhuXPZhO5dV4QQ8nUD
eX5zMwgmKbhXtQrwUW3oBWcBekyA7iNeY2dSlRkzUIAAuwCjaXT39JcTC8vZ55/2xjo0Mna+pC8+
7bxosMzUIxsZbLJ7y8voexky+aOmFJn3RUzFJJqpm9SeymiAObvJx5QYaKc1oIpzRgzLqPtlr7q5
fScr1l9a4GlTr2B6mj4VRQtKAOBYFib0IfbsICkN/nP6mdHNj6SvpzwZk4xylHDhaKYjdf7cpjvt
ZZeSqQZlymxWyXjeQz4F3toaXQx8iQNUNGCHgKv6NuInjbA4NZ0rpe+XES9tLx9safQVn4IPoHtv
BWNLOh5/j1xFt/9P9NknuF5BNdy3EGwmbKEFCZoD05x9uB180lGO8oE0Xk9hmYPjFWs1yeZiI2Wr
N1YEPCUXjyjE2Mxm65I6Z4lESJKIM/aRml8ZQ+dSTMe/D+FE3mi7ksRGinemoYQU+EIUDyuZOR2X
djeZXhg5kOcWtxtliI9PFJRk6G2maAKBY18EF+HCy7DyQId/6gOKa+pQHc/yhiRCcEHRf4b6A6PM
qZUpzoRR9qSu3TsHToxXRFx70vL4ENHCIdYK062veBPMeNWb83hqhDoyEf25l5+462y35MBvJsE/
j4fl7ODOS8XEV851bmDUV/OSQjb5N/sp5cSRAT/13lXFZY/9jeHdgb5bPhO8mYGLn2oAfldPTAVb
xO2BoHStROxRciNveVRjyn8p0aE6UO1I+AI8MUl6xwkHCbda5Dubv65EbA7ld+/loA6TjLNGzgLi
pmuHFMldWf1jWZ3oFbHzpKmCFtwj1+WLd3jggs4u+hJlIEMDkHjAfzfw9g/tNf4t4z+lFuo6InsH
clmVIpFVO27IDy3k23Xsj96YwOqpiE647V7ci/ldph+TxtVHnI3V8Y2sG4vtn5HmPmvPrqhaNbHg
mY1t4BMGfzhbXMt1DxxQoKn8J8J/TVtOhl21e1Wcxf2cmltkVzoLBm5pKlHtqJkRMiV+mD6ctpY0
89vNGrnbXMTzQMQcE3RYxfXQhURwuhJufQaMMu7kC5gOd4nBz4C0xqcqFHn1aNVipRrzDm7O6A0H
uy6pDvXGKdmDN+WRvGOHMAdzBDls+ngNtxjH8mITPA60j/TOTgpo/7+YSK0eYAUQ43suVRtaoFxq
Wzd2QgvD1hpRzZvwA7Dn5E1KmOMbYsB6klECSI53yayTa1fzZwstxoDHf0ozNu27gWA1RGgPGZOb
7vj3McmvV1J/tAsj1vKaBsZseg/64kAYyqD2U4HaOy/jSQHN2ve4+yWhs0Vcc4ZVltBnmFaxiQOV
reSjI+CE0QQWCwEzyEJPERZgPFToXm0Dt8Sl7JDoNCG4wG7Fz+E1v798NqE2uj9qt82helxSYzxl
Zo6uuhufaOY00FdKVUCsLuU6KeUmEuhejdIDhDMZ5WFLHIbFiztfJ4RGbWA54F8VGoZaDVk8zz9P
/A/nLZ3KsYvZfcICkZ/ryGYvRIenjXdkjei32IS7SIlreHmLwvTW0l5csnnWvWgqtTmdlpFcYOcb
MQhCJcaDP91hofuqb5cEMTjV4gwys1GG2dFVqdY63RnmHLm5gEFnAks6ksKyJr1D/Ttf4bb1usd2
L0lr5O7DdpLtDAQ3sBuXFYlJ8xD2yfvM5g3CEzMfheBIhAHOWf5P0VlSU7HZ5gaQO+CIScU9jruZ
9HZuX2EbC8P0fYMXQsatTdRRXrRDQIEffi/9w6ekWLhlrHi7Qx61H1T5+cQpthllLYIiZNwOL9uM
ObQvsSMWvJ62NKnyiMylBuTtpz6n2feYZlyXonrNVbttVkPiqW5gNNrZGpbnO8BZ2kK3UwFf1xfT
F+mA485z/FINh2h2q2s8GMxRuQiY1o0PrWKtTUopbjd3ujvsuTRrleCPYvVe54GolL/LJv0XWTRx
cJlgfUG/vklJj1BfdC7BAZKz+/ikfOD9FLTNlesm7GJL7BFvw/96g9nqAJAHemVpihLi9W4btL6F
iAhFbHIBr9P6ZxiPOnLeFCyAXE30j2uuCpFfAP1WicyjrpNqmne75Wpas/NIx8snRycJ95svdH+7
zt2PCKceftR8plir/EZNVgKiE4dDQHeaRcOe5X0ZXQBzRCfjzaDlb3Hs5ibz6L+duNA7AXexe15W
rvVioDJ03dh6i+JT/4mHCFtL8FwXIrkVx0rEz98t/9st9NpNHy/kFi3yuF7zjltKzCHfvVarisr4
pW4Vt4/gmNPmvs7ozI0bjzzBoRz3S1DkPBDHdg5McCJKlaLcfdjcRqB82Yuv0OjKY14jfBLoTAqJ
RUFAREKs9ldKWXzZgWtw5kRvuF9ceYYEvN8YKtklJHNcR12KH4qMNWi8TnLdZKKOzEVbYv26fb7M
nHoyGv1rFturOLxkX16PgciNP2qXu2qX2UUWLnWRb110huVGrdzahWrKOX20yiOLstKLSiHewpTL
lhkoJZ1oWnkn70wDUe8es/Ib09C732oYUL/HCazWZyF5KtPOAr117HUQZMgr8HaJYC5LeBSVd9gs
RPtv9Y/+HZ1UXixswak9dmiNCC+SprUXzJlLBiG1dP0gvaVTwPOuxRH/+sLrjVJ1vdCGA++j7O3Q
J330087I90RNATvSh9czctOliJvVCudCCMvIf/aZ1QO+qTIt6mYSqoxH3t+vHz0dKiE4AFZ8naiq
0F/0OONnUdbCOQU4DpdiJa87pVCMrGPKE7w13vRRcG9n2A6p79U67pKfHPBknk9huezPrKE4qqkF
HltwOLeQ7wB+iJhikfrW6NyX1lLJyOTnicnFeYIgSmkoa8KW61sfgazybFNc0L6tQT3dIOcPC/kx
rMJdBBI2c9Bd4pyh/nCpWx/r9/DKIOSdYOkVWYZ8ZyIOMLDrzvuNTFX96dKm4kxqCgwb3vHXYHMP
Va933iGG+a5P056qSHwpinp1Qvth/SR9JLqPQ1KPXhaKF22e3RaYEEDHX1AS5i/MFoUBXL/3BrQ8
aSgTZQhgAWhVInsV9tqEaw/mCs+o47DunQXSqSlo5wwA+ASXQWT3QPJnuyrRih9VOWr9mNMU+iKK
iMT/60n3uofqJ4GRchLQXEHxIMlE1i9MtyrLeO9yWuegxi1rS44X0ETQnOmyxqhPYPTLIKHFc8bN
ZG1Wol66sFXMeDTJ58E58aydXCNVJu3zH/RY6OvvOfG8+mMyVjzaDZhfbiwU9SDfz8DwAT7IroW5
DsqV9JwvhdAYU25QrkXSehjUOHkIU6PV2a4kURnQZg4efgQ9Z7LWdiTPE4laChGCbKJr5mpHV60d
tN8eYIOq8TmYhkcMju0ANS2wxegywyHxaKGs+26F043fhUnss0tvw4k3I0oYUB1+vgc6/MOIN04E
YtlG2RxehvE5oUvIc0TX2k4bQ3NVqUWs2oL4QARk6+EWwXb2Qecwzu2FHlGm974E+cO+bTXtvqa8
r45pdvOPXkkgg9t6J9/zIXJLgP5zjHHQqT0rcBr/kpSwhIXdDTT/0oKBe6G86DTaptL5tyTEEPKS
POdYB53ysGNFpy+Md6/55ikiwqSQKj/arsoj6MHGk2XonUOYcW8R7f19cm9Vpc5L7JtCLD/3YCGb
+UkYCh3mYDhbJ3I/RdtVUiIh/5L672Vjh5yiLyb5i+MtKFyIPu4mOd2N+YYDe3hAl/qkoe6OaYcX
i3H1p12Z3LXKIsP4IxUgwZYQ+4N+wG9N538lbrbhyzpCN9wrloEz263p14FUemLpJi4qfNibobi8
C+WIjlJ4KUexV/UJixq3hywcaU3FEgHnQLot500EXh0ig9Fr+qwyREiWmPYb9jx6OZNFbowFRbml
2TvNc3xq/4skuXq7B3cilb5UHhbvycq/iZF+azoat/f3cRrBN9iNZ/7sdlIcVE8Ppjn1YRrh2Th3
HoAqvsr5sEA1LUlhMWjnW5zPgYwgHdGjyW6s1C4Clz5lU79kTwraARNQQG+FtXljsfDwch7x4QMV
c/tBhzMnpzKLUWWW7fiAkGinX3qriOqKACujqbdh8sZRgumTyRLnnW71S2faIXBsgmLkGkrtxdxp
CZUmRjXKx3pVoQibmcoIPfEOXN9udnjCdh+O0pEZzYzzjPSqWP6hWIwkZOYNQBjM8wZPqWp3J4p4
u4e/62c42xMtcp5xgxJH5ykukoY/jmBhKM8SWqEelQISQfsBNPXZRoGmK2aw9p5XCyNUb/C80h0Q
3Y2hGSx+y3ovvvx25yKx+Ju1funInJiFCz5whwxX6TcKDj0XnwOEbmQs86G2mNTD/vmA9WscjqA7
/NjvWroGQPh6caLEX5/wwA3jlwSX5vn6yfP5q6r8jobjxe2b3+Cwg+qTvTxyc0yDXxKbGw6TIcFZ
N83iph8WzkczfO4EFDLDc5a6ELcqULlD95ZuZdsnu9MLboEAfpi+B/s6cRaW0uVmukFhEaHUJ8EM
xD7qFfqXz4eHlc0upjrOZjN0Ur96yFkiu1rCU5gnaYWH9fBeiGx8EI4WV4P/9QmiazD8jNoikNzv
4xQ3OzRZ9N4XnO9amwBPxth60y7arpyPwqK2i4yudSERWNPb7B2c6J7k/Ow06kwDrIxI9X5CmQNq
bFzYdV6lHxL8p9/mRaKxMkVB6TBADE0bAQoaQnOZHooOQCRKJ/v32Q+1CYsVGtlZjtsL5sPaSSbn
L7UdfmGkOBkbXP7S/V9GAhTTQYxoNzVf5+tIu6b12PV56hQohC4GKUrHvFujEAXK/Bz+u+LpWOYM
EgJ/pPwzzNtnXwHpW4gUi5hHswnWqv6XLwyT3F0wznZponO8H9rFkczc3htpUrsxBLj3t2F+bGbv
M6ONZug2qBfVwd7Mx3ZQcZn2Mc7JWKd9AaTCVJidyzft98RV3iqU6ibQTOj3NAGJBqi35jg/L4cf
i59BIO+ba2eAlzNc4Wg6UgHnLQrEOXeQzT87M8gsrc8k1qMDU2XBT/LrmErTEj5KLqV37HaRa9U9
H5YFM4JQdbY5ML3vfBltAdyOCMeq5TNKrFNYytSqCQd+dmZwERpbmv+ydHjyUtAeqz1hI5bmcCem
xUsmPep89BfEoaThmMM3c6unDsHItQ1063A/vdnxYtWLa7hazOtjHVERStlzIW2PZVwPAehLwxgJ
H1lw30VPTXFD2sKKvdlB8fNykaZZIOvl/1YJVcd8NIajObkftqHH0Up7G7MaAES4JT/ZxTb12Cg/
zhzSXW+tPvR6/p8rtidyd96j6m3DeUPk+PNfzA+DrDtr+g4nORQEnBpxE+/9Vzh2urDjY8PegmDM
GUEShEoIJiOT/yYpaj8g5ZeRkEURd1hWLf+GdrJVmayDNpGb1Pye2pzRd/AWExlRnJ9XQ40L1lUg
HRv4Ih5Hjdp3q10bHnJQrdl1IRLOPjDb9oyvC/wKB2sBxS7ObMmdKj7b/SlaPp17k2JavPmOBZj9
89rHnFqifgCa9SpBXwOM3eL5L/AeQl+XR6oE6ULGRgMdmrchCEaoeKEP8jIRsJF569bLv3qcARvn
I+u1phwYjgKrroR7ARAvGWO4XK/TEbPX+WKwI0F2Ba4D2BnetXUUp5howco9f7ALO3JOF9d0K+xD
NUOeKHSQbdEfyLRAcm3dlfKz5TzHolti2mGZFRB3TCy6YAm8Ki78zy+XT3GRGFEROngapf2KYWOv
V1r/bLV7FiNVqkIKx2ZlRE+rTsNhTtjVjkmoL7NkMP0eZEYTaKXw0eOGDu6zNJKdk8VCqDnMFhjw
79PNd6MC8ZBU7URA8eb9vRekD2YXHa+M45tYKuQAk8RAahSp9qK0hg7k3iTvpkWRgWJOo7zTBDnR
hAsIxq/xZlrlDuXGNtM8JgRSkusuBnPDnyin6xq1qewxtzO4nWm2iS2YICPP+HsCw7fhFmMzg0W5
NbBjk6/g9ueBANwf63/ecQZG43zergJDa1hMRZEgz381KhxvZo1vsWzTY/5eq8+BLlTtR3IwZhzi
ydYLO5zqW80ahwUoq0yiTthjfaAki6pGWZpsDIKnxO+lXTtBYxErwfKr96S8RBYwA6xUuWMT6rzo
PmXLmCrjEzIGBtefiR18jyNuDzBEAfzhwJCx6XOABJf6kOXnw92SOOLt+TKz0em64cQ4ho2opR+t
GdpOhJLrOm9ERlIsUzoKrxr+pVv+IoExtwos4DNN/X+jnLmHxeh2Cg/m6feu8gX6k8w1m7L8lWFI
+A2pgUkC9x1fPaN7xzLcqauW/da7svw3boJlz9Hrgc6WDz+DgmRY92LWcYWLrgXM3tjZ08n5fMNr
WR7VqjYG5yIEwyzwokKD9pBc4ITuKDOwbV6OQSyKYVaOo0X1ZnEqKLCVjixeME5QZAwKiPBOIISB
u51bySFI+fQYGly+3BDkXmgBuilUmL0IJXJ+bFDFCU+orlnBOrss9CwHupiUpqSeEojB8dDO+cgn
cIsH7v0VYX3vZhdsQEj0zz0I9VINYO0NDi1ykU9sGN4tm7LvzQ03WVAHs4rl/E6XhilQQZi5qK/Y
J550AbrmWb6UCIOVqySw1ZwXn9Ex1Maamvl5lgTJEpN6wmH0Zb1F
`protect end_protected

