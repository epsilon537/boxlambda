//
//  A simulator top-level wrapping around ibex_soc, instantiating SimJTAG.
//
module sim_main #(
	parameter int unsigned OPENOCD_PORT = 9999
	) (
    input logic      clk_100,
	input logic      clk_50,
	input logic      clk_6,
    input logic      rst_ni,
	// usb_device leds
	output wire        ledg_1,
	output wire        ledr_1,
	output wire        ledg_2,
	output wire        ledr_2,
	// // VGA interface
	output wire  [3:0] vga_r,       
	output wire  [3:0] vga_g,       
	output wire  [3:0] vga_b,       
	output wire        vga_hsync,   
	output wire        vga_vsync,
	// SDSPI interface
  	output wire  sdspi_cs_n, 
  	output wire  sdspi_sck, 
  	output wire  sdspi_mosi,
	input  wire	 sdspi_miso, 
  	input  wire  sdspi_card_detect,
	// Audio interface
	output wire       audio_out,
	output wire       audio_gain,
	output wire       audio_shutdown_n,
	output wire [15:0] pcm_out,
	output wire acc1_overflow,
    output wire acc2_overflow,
	input wire 	     uart_rx,
    output wire      uart_tx,  
	inout wire [7:0] gpio0,
    inout wire [3:0] gpio1
    );
   
   reg usb1_dm_host_i; 
   reg usb1_dp_host_i;
   
   reg usb1_dm_device_i; 
   reg usb1_dp_device_i;
   
   reg usb2_dm_host_i; 
   reg usb2_dp_host_i;
   
   reg usb2_dm_device_i; 
   reg usb2_dp_device_i;
   
   reg usb1_dm_host_o; 
   reg usb1_dp_host_o;
   reg usb1_oe_host;

   reg usb1_dm_device_o; 
   reg usb1_dp_device_o;
   reg usb1_oe_device;
   
   reg usb2_dm_host_o; 
   reg usb2_dp_host_o;
   reg usb2_oe_host;

   reg usb2_dm_device_o; 
   reg usb2_dp_device_o;
   reg usb2_oe_device;

   // jtag openocd bridge signals
   logic 	     sim_jtag_tck;
   logic 	     sim_jtag_tms;
   logic 	     sim_jtag_tdi;
   logic 	     sim_jtag_trstn;
   logic 	     sim_jtag_tdo;
   logic [31:0]  sim_jtag_exit;
   
   SimJTAG  #(
              .TICK_DELAY (1),
              .PORT(OPENOCD_PORT)
	      ) simJTAG_inst(
			     .clock                ( clk_100              ),
			     .reset                ( ~rst_ni              ),
			     .enable               ( 1'b1                 ),
			     .init_done            ( rst_ni               ),
			     .jtag_TCK             ( sim_jtag_tck         ),
			     .jtag_TMS             ( sim_jtag_tms         ),
			     .jtag_TDI             ( sim_jtag_tdi         ),
			     .jtag_TRSTn           ( sim_jtag_trstn       ),
			     .jtag_TDO_data        ( sim_jtag_tdo         ),
			     .jtag_TDO_driven      ( 1'b1                 ),
			     .exit                 ( sim_jtag_exit        )
			     );

   always_comb begin
	 case ({usb1_oe_host, usb1_oe_device})
	 2'b00: begin
	  	usb1_dp_host_i = 1'b0;
	  	usb1_dm_host_i = 1'b1;
	  	usb1_dp_device_i = 1'b0;
	  	usb1_dm_device_i = 1'b1;
	 end
	 2'b01: begin
		usb1_dp_host_i = usb1_dp_device_o;
	  	usb1_dm_host_i = usb1_dm_device_o;
		usb1_dp_device_i = 1'b0;
	  	usb1_dm_device_i = 1'b1;
	 end
	 2'b10: begin
		usb1_dp_host_i = 1'b0;
	  	usb1_dm_host_i = 1'b1;
		usb1_dp_device_i = usb1_dp_host_o;
	  	usb1_dm_device_i = usb1_dm_host_o;
	 end
	 2'b11: begin
	 	$display("USB1 output enable conflict");
		usb1_dp_host_i = usb1_dp_device_o;
	  	usb1_dm_host_i = usb1_dm_device_o;
		usb1_dp_device_i = usb1_dp_host_o;
	  	usb1_dm_device_i = usb1_dm_host_o;
	 end
	 endcase
   end

   always_comb begin
	 case ({usb2_oe_host, usb2_oe_device})
	 2'b00: begin
	  	usb2_dp_host_i = 1'b0;
	  	usb2_dm_host_i = 1'b1;
	  	usb2_dp_device_i = 1'b0;
	  	usb2_dm_device_i = 1'b1;
	 end
	 2'b01: begin
		usb2_dp_host_i = usb2_dp_device_o;
	  	usb2_dm_host_i = usb2_dm_device_o;
		usb2_dp_device_i = 1'b0;
	  	usb2_dm_device_i = 1'b1;
	 end
	 2'b10: begin
		usb2_dp_host_i = 1'b0;
	  	usb2_dm_host_i = 1'b1;
		usb2_dp_device_i = usb2_dp_host_o;
	  	usb2_dm_device_i = usb2_dm_host_o;
	 end
	 2'b11: begin
	 	$display("usb2 output enable conflict");
		usb2_dp_host_i = usb2_dp_device_o;
	  	usb2_dm_host_i = usb2_dm_device_o;
		usb2_dp_device_i = usb2_dp_host_o;
	  	usb2_dm_device_i = usb2_dm_host_o;
	 end
	 endcase
   end

   top_usb_device #(.J1_ROM_INIT_FILE("j1_mouse.hex")) usb_device_1 (
	.clk(clk_50),
	.usb_clk(clk_6),
	.reset_in_n(rst_ni),
	.dm_i(usb1_dm_device_i),
	.dp_i(usb1_dp_device_i),
	.dm_o(usb1_dm_device_o),
	.dp_o(usb1_dp_device_o),
	.usb_oe(usb1_oe_device),
	.ledg(ledg_1),
	.ledr(ledr_1));
   
   top_usb_device #(.J1_ROM_INIT_FILE("j1_keyboard.hex")) usb_device_2 (
	.clk(clk_50),
	.usb_clk(clk_6),
	.reset_in_n(rst_ni),
	.dm_i(usb2_dm_device_i),
	.dp_i(usb2_dp_device_i),
	.dm_o(usb2_dm_device_o),
	.dp_o(usb2_dp_device_o),
	.usb_oe(usb2_oe_device),
	.ledg(ledg_2),
	.ledr(ledr_2));

   top dut (
		.ext_clk_100(clk_100),
		.ext_rst_n(rst_ni),
		.tck(sim_jtag_tck),
		.trst_n(sim_jtag_trstn),
		.tms(sim_jtag_tms),
		.tdi(sim_jtag_tdi),
		.tdo(sim_jtag_tdo),
		.pll_locked_led(),
		.init_done_led(),
		.init_err_led(),
		// VGA interface
		.vga_r(vga_r),       
		.vga_g(vga_g),       
		.vga_b(vga_b),       
		.vga_hsync(vga_hsync),   
		.vga_vsync(vga_vsync),		 
		// SDSPI interface
		.sdspi_cs_n(sdspi_cs_n), 
		.sdspi_sck(sdspi_sck), 
		.sdspi_mosi(sdspi_mosi),
		.sdspi_miso(sdspi_miso), 
		.sdspi_card_detect_n(~sdspi_card_detect),

		// UART and GPIO
		.uart_rx(uart_rx),
		.uart_tx(uart_tx),
		.gpio0(gpio0),
		.gpio1(gpio1),		 

		.usb1_dm_i(usb1_dm_host_i), 
  		.usb1_dp_i(usb1_dp_host_i),
		.usb1_dm_o(usb1_dm_host_o), 
  		.usb1_dp_o(usb1_dp_host_o),
		.usb1_oe(usb1_oe_host),
  		.usb2_dm_i(usb2_dm_host_i), 
  		.usb2_dp_i(usb2_dp_host_i),
		.usb2_dm_o(usb2_dm_host_o), 
  		.usb2_dp_o(usb2_dp_host_o),
		.usb2_oe(usb2_oe_host),
		 
		// ym2149 interface
		.audio_out(audio_out),
  		.audio_gain(audio_gain),
  		.audio_shutdown_n(audio_shutdown_n),
  		.pcm_out(pcm_out),
		.acc1_overflow(acc1_overflow),
		.acc2_overflow(acc2_overflow)
		);
   
   always_comb begin : jtag_exit_handler
      if (|sim_jtag_exit)
        $finish(2); // print stats too
   end
endmodule
