`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LWYKVG8dfc8ZspadWNBtxbVJ29EyboKS0TaMenpX0CY4ADyQRo4CzaqWyi3ctiKvT8t6iAIl8vry
qUuVkOJL2UhQ4LKGDRgQowBoG+VT4ZeQ5JY53a7otVg1Pa5Gy0QanS1PTWAenp5vpggn5Tv5N29R
Ok62KfQ/E/p7qBO8DKF8s1K5p7Sf+tGAoLZoSrU+y9AzQ5Red1v8vHy1IW7ISAGKrdDGrK8siXq8
VVR7wk/kCjB6gneeavi2mB/R7TNxoNDeXxAh397hTfwJI3s8Mm/nr67HCyXJvMDw9pgU5U5s1Kaj
GeU9A7iow9cyOwYQ4pbqH64A+CNt0NXR2FFyfg==
`protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`protect key_block
Kj/SUF0SZZ9r3ZVlt4BBDoloHfwWWTOK7L2TkVUDJUQsn5qe1DgbDGk1pJ5QHVc8N4/HRHrkDmSk
jA/YUvDhAXOjmAc6DEo1CtJkT8ZlBh4yns4iby6hiyNCZLBKoZ+dc6E1bcPOSt8QG5d+doe8DL7N
fjV1hfieTn8Czn/j+9evtsNeqG2ttx9NMIb6IhUE0Q3YXimVuYCcrydE9Dvi0KkMwFC1OCsrokPx
sQEPShPMx/GHLIwUblfiktEIloybb8HD5qCo/55qlj5Z4p3x0hKJ+LhA+jf0aU+lWbQOED5snobO
qZRE2sd1FoANN9Q9ttmc8742qoqIidGvP4JavgAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
i1DoJdoYFCWmKOq9GgqeHkiyxL44IMKjlFcVZf8c47izrQEZC1b9lsB5UYLiNSiLlJA8Q3tNhYou
C/QidAcweA==
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mbPfseFlHOwXfgkW9W0yIsH37mP52mZUX/NiCZd6keezrXoEylRYINwbHmdtk97MO4/YDSAdLvoq
rx6FYH7ibpm8msK1t3PlCLIIY8ty4+R35SCd6MkfudqmFWIJ/GdrofoYNyRsR+fqfws+E83rODFn
AnvsscoQf1HyoNOuyiKlfPULmlm6ZO09rLrMEpBWhtyxVaVfjaPMAagwNE8boRmRdtTjdjTFrYiX
lmC5ydT+J/3pbYkKLXcNtc//cI3f6AtbVz6pVfqu6gvGrfNWByScO0ByUW6DSdlrQtQU34itPL/i
fi4LmJwYcMduUaNX8U/SAi/BDfoBqGJ6ER+FBA==
`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ip91dsrln+U/dZr3NLK0GXe3y4pWO3NRb9SOs9abU9QBJa7rAxbxOAuzvG9dg7QvKcdcIlik51A2
rQ6T1P66v0RtBVmuUBU/3uZRcRN7Ce6QZ+niTko3tTadYWzP/BD/wssihTGTo11ofvKkpTS4LnJ0
KoDsGgbFqoQUhDHomDh39qQm1wKH0AGvVuetyE80prpLU+Bi79i5va7+YFHNQzNJ9+bqh8JReRHB
COKDaAg6GsCgo1H5KDJLJD9Q4tfKD+i2GXyhZmAxHgFT9p3I44Burv+JFXv3OrRfdA8S5GLRG4Um
wfs2jkjLaikHNHP4gplZpf8hG59ia8Nb2JmMhA==
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
shCpR9B9uP9ZkDWBHeccZL+6vxucMjGwubE6xyHiGWQSGEy1q3KO1/t9gX9CCT3dhlF99CcSj2HW
VvDv6KeFib/+64CZJdTKhQxabQ49PrkOWg26TKTkZkmtpfNL4g2FP+ghZ8SaLeT3FgSKNauJqPDh
Yu5LQGhqBCQSiZ0ZwZk=
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fnnWxjjOYOFmoV71hJ80gwYpRuTOHH9EgeeKMg8rlcHN2EUdpdOnOAjKLqHheBgZeAWrz9J6viQa
zEjOhgMCr5lwxbFyVc70r7AiU4UuaWbgkC0QyEP4EYOAY4ADHl/9YwNv1NdqLx6AKhvxkchqjgqx
WcUwj1IuZt3gJq9BV378Mna+yKOjB1Fu1Rcce8ChhR7YG5wsGg4zrtgoTFlYdFUoBpGtgWtNHLy2
7sV/FuNzqhSKdagnvIZ2D2vEVYquiwAKybMC0f5D6Y0MRjeQjU/WP3awJRc7/0g78hV1wrzW0D/q
yyVXeCObqtbXLSuzj4oml3+zZpv+Nk+cihVTGg==
`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Uq+JLja7j7zrfLbVXtpNfPDm/LASxfNbBMlz5mkHQNqBpEO0KslIl2rkDM9FHXn++FXAdlJLhg1C
et5vf1Xbjh4XAvoNStdf0zDr3imK4bjtPkMDaCNGbc+NS1ou2JAOnEMVF3RQ3jObo7XIII/m+Snc
pQme5L4rI0WgyBLODf5GqAfPXMPl/SlWyKkk9k0iy/N/u9v1Cfnn8O3+hnbHGST5Gqgq8joqErvF
qusW+PFPJ+5HgoByPiqYAioM69X2fDNEtzPNTVetDLByoq8wlGfdVVi2GAGj9/ldDA6cb46Dke6N
O8T3Z3PUOQ/h7QJgw7RsIFIeMi7mSjR1FkJbxw==
`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pZLTqOPhpeX5czPwqf8PqB8uyLRrnQkxtHYlZv/vJcP5oQc2EWKcbfCYc7ZmoWRe6xIW3kvT20cy
jNVzTnnbfjFXX6aIDfnl8Z/0Xe9ymBR7qEwXY60Qx5JtTCVlrzcc6wBXGBPRTb9gPIRcMnwEdl+i
/vU96U0JTm2moWzBDbI=
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jsxwPnal+isiQ+Gf3A1++FQeJh0heEVAjxVGr1+RZQdUWHFa6pfiqLAfbGb+yq5/t2ruz37jgntg
oCZ0eXsNxA5oNwcC743bdbVCbv53WjMsbitjduvMTTbjpnq9e2A4SLC/lWZTJX25VLGSXVi3btTU
O8YA2OmI9NUVaiqq/Z2g7LtnJ6eHABGniPP7eyaA8BUO3gQbDrlDX+vJNinMFDzhjzLTDEHWbb1B
7kHT3VZMjxh4xpXCHTivHiCXKdOyr2Zk8rv5AAiU/YJniRzYB9m8o1/jlYPd6m620AuJl7O1xr/G
QFUSFuDFZJzMuU2F9fSYNhoQXCqAxK5MV91bPg==
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11888)
`protect data_block
4s2WZZ0Wf6kwAG94T+xYxa3YU+v5qzKxKbSIskcL4CsSObA+pHpziwcuIs3/v79s14MO1ONAIdlY
FPCKNUEpd7yD1ycZVgqDHEUVY2X0Hkfi01zBoGnhM2L2Wxo0VWd+mR6pOi8KQ2ZKegQZfR/4RlLY
8JwMhI2XbE8HT/WdM9E4zzWZn2kxLVV16LavcPDlgBt2YRQlIFAuwwmJRxSMdEeiRNAkV0vrHoEK
K+Ijnob+hV7ZkkuNuDymHEWlveZpR+VZrkxjl4ovZOMhfvhHpmrwIb4tx6vr6s+NMlJErR+yO5/G
pLyZTBlRQcHK9PZB5x7jEPbVejFwvVfbXRwCDncZnHXhBnenoU4KZCi2Umb7ukXVCo11uTcfZ5Ey
0bxKmSHzGRytSp9GrM6spa/7FsryOtLyxl5a9l7Z/Cy6k/jqVn3L7PkalFmVR+DKNWozRhErcIln
FHybi5MNDki590Pc0MIwYXN6BrhL2beQwN9P0Fwivjq3GpgIrrw0Jir3J+SBcB0oPbrxewl2QPfO
Rnuvq+wy+lNGrgpG5tgfbPiCyIVB63DjKtkBnn1UU5i7Qk7SlIjLqVr5UKM95/HRqKS8IoSy1Zf9
GVfjsIB8lsVgoAVSRVw3d+gIlE0R9s0NshWyH36tLbNkclCM4iJFOKgZUEhOYfgszi+4US0wSuRi
VQYvuOAHMwyiIc4DFPQOywsKvW7jwahu54bDS9svTW7RImGlmZnkQP/mVuXdMi6xVopnmD7Ixq8v
/Wxrdl52C9DnfN9uW7f0Xc1KfJct1RhgEIWHmpFQVxE0It3SqeUHpnfzcwFtu+YT9ftOjW78D8j7
V7dpTzot+kvVRAjfqySIAUwj2+Dik5/YfAh7QivkYzeFWOpeysizTJsEgxvGhRwZEO/fVMe3kbp4
a9pTbAJ6xIqdXMwlTKlXCYnOFfBLTVd4cUiybAASWYu4Fq2dYCB0zNA3bn4w0GuujzM1b35cvhgi
apF1t0v6iVgAvxSU91ouf/cPPhv22zaBshlDlZg0TDA+DTCunUPOfUPc3tPxWCJiO0f/NCXpYeVb
58q/UjdznST0MGb6L6cCMwN/kyDpDFJFEyaR+APAnAJ025enVFX3Sf7JdWQOu/TJOZr2USyVDBtM
IIVqh7N5ml7IQkVVk7btzv6kzYAC7lC9yEHV1ekerCDocP0CYL76QC1FKwsLVFcxTuuGYrWqg9yC
e+AbG6uWpLr+GYL5r1RBzj44M6WLQBvPdcNoinZQxhG6aDRxQX0wF6fHCLYUC1KyIkk+rFv5BBYD
tJDaIX1l94I3TSMNeBUjalytkv40eEFWbncvg0CX1Ut7OWGrIdwEFI0AKQ6aQ9v2xfdkLh6ht6gY
rHY8Z60z2sHxBDy0Z8HrqMX8jctKJudSIgk3StYXSTJzG1W+b7d9nmu2gkEvtxix8EEAZuzDNVQd
EQ9y1ZWTn/jShaEAEbLNXN1qSx/dHSE44VEP65sg+T0Vl/0XbcJrA/MPJ0G39E2jQQHd4d5POPAp
aWk5hgn7deCDx/9pVhmC0i8ZXnq6LGBDO7Ye3xFZLcsJbLyn6pbMGS/HcCWAurax+pCqSWBC24M6
Xt3hTrFp+6jS9ayVl9OKDOFJdPe1nrvpOs7VMAOyYBxLr49HMSUSkqk7C32XSv3mcp28Fc4QfNrq
HLUQTHcWzSLXj/8g6O5GKxfn0Ef8ZZ3Z44mz8OFfOZqMEYCYtAwplWNCex7BAbuV2TsbZ/lxwn59
O+Hs0C3vHVYC8p1YkcmaTwEXkVowkhfKhTgg1JpWynxlmiYeBfp4Jerc6AK56//45cIJ6vpQHo5V
G861mW95pq+Bv0eUvbCrHJysgNgysWa3M2fcy/pieK2r0Bpsqkuah0ZT3Jb6iIfQbdYjMWCSnVuq
+50uq2cA7FuDk7JzHaCT2uJJd5MuBO5jJAt41r7MXnIBWc91wBufkiIc7DgTZzNO3KW6o9j5LSo7
yTIWQsewt+gKsdkbQ/qYcRg8JMbozX7QhUsMeSEwJUNDsOPCzc6h3NblQDypjR7zZkijQu5R0444
lDL0AJ/kjCG5nbSAtKZjyF3bMAAPPqrvsMO2zce5wUgNVmgRrsGZupJTsxrkBcZyWEsCiA7LWqpN
bK1+Il9h6rAaJT+kZX6OITB8uMFvKQd7XAqLzaWeK/hyzBpTAwk8DGJOHnPX2hhRM6CFEktr3WJp
1ojwOLVqNk9wpItlo0zccPjWbjeRFFEWv8FYVDbiAQLNfOQUgbPWUbilhuAKwIMeaDNR2Ir8HL1w
vNb4xgfRdRxpnfhftfnIUOX9y9+bCuTSxa9z40bmZ875v0QkmhPKohGmfoG90hkI2HicdDu9oDBZ
iQ/eimZLlIl6lnPzjES1WkshtqUhlEz/iCViYyjP4Sr0rRhEIZs9CmVjNWRNYFkgWk8h6TALBdQa
zDxRkJcWTRj6b9rPXIUHi95QX8vLA7cw2CvJXdd8fBcFk4mrsihNGIWywhT0J8cd14BIWE1jk+qL
bqfP0Jy4SCSnRf3OlageFacgtYBLQY0VpN587JNEtBgBneQ6z/qacj+ZnGQ2yM88m/ypxRuImUD+
LQFAPx+3PxhBQRlbEx5Ls0l7sds6InpPWlYgtiXcCuOVYTf52Atn+atmmolAkDD1N8MiLtjRE55d
cO9hPAhZ3PT54xTZfdGVr1RebEnrc1/2wVYfpROdn1cag91EidQAQVgaRN+6qSJ+3h6lpYJR8fPx
XPzdrZDSWwAe79oq2aGO+0l3uKagkuwTZWvEfI6XGvEKKhpc0XaqpTfPL8VI6WFagWjVjA1hl5DG
bVQRrEP7IUeJ2ISFtqUh8hGjgj9PP+Tq7w3AHABMONU8caiRN8gnHlzF0ap/qvEMruGTZiI8DHVo
qZ0MMJ1CNJq8LoJq30o5UY1L61cyXhegqbxFuHjALrfO4WjBzscCVYsHEsZ/2g0dEXXOX/k94Vzw
JxYSp5Lho2KupxOOF1bhavUykrAnjCqUWUvLmXNYJW/5KkTDf7oXYK1Kp9PRpRRxBCG2Pj8F027l
MFNQvlB8F9hBk90rHDgbsopcWszsONdmVg2FwiAgEYR/5FkJJ/Au22tE15ITuZUuLQnWySxqTHtc
mOBZ9q/tvRtc3ZGQ+FUhG93FD1i0jvYg57FNgFDk7giOQLte+HznyjMI+D4cDetUUsrqupwvofZh
FUW+58SYsGBa+aQuF6vplYzL+ASre0O6dJvDFZqLZgB1AuiH7vGSKuq+EuRf32NPRLlLI8RltQlo
eNrIA9BspI+kMfUdeEL+IlIEdZJ0lqX7wU8Wllk3FBS77lkgNy5qltyzFnvWSKOZqV8HKC8lGDdS
wt+/m8Ps4BnxGEXDLKINGRKkYemS5xfrptYqeYqcJp4xYT7VVGiIoircodGwnq6PJlwpYNtMliag
oBWAIKjt5t46lwqRW2M9qCHQaOdzwQ8+1emhF5rrZq7FTQ4mFzMdls1Nkrl4sPoYI+A8YRGy+ybM
HilOEdniWi5dYH7bhAcGZm8/a6knapvH9tRrsoNnSPCkZxJd+nnbW2gpC3+FpmXsaBotnwdZRQWD
uGzug1tB782rpAjdGbB9sYj8A+gU10NPCGlzRilHoYC7ut7HGJfKAN5rISSYaF961tBK2VuAT35s
rGO9JyK1RACUxOsyh4J2zkBLzup90WelkR/FDcCFdWR7rl9mwmMtx8DdeAgHHZwnkL+AdZ0Gi2Hb
UjdF22myAHpw6LLzasQMuoX9IKG9NemTCHt6me3Cakbn8naCzhBU0iGfdZE+IbHtlJAwe4vBx4IY
4nX+EUIwmSjk0edVxSCBXbh1SdsR4qwUUyBoj8psojgZAzYSh841SHlfk6k8x9yXthmwMdeAU1FA
NhSpky+VvSLCj+Z6vBdCn7aXOIBKaVziTxJe0Dd/uZ09li2N39qo68epdT3aEminPOrPC22it2gd
XMXQ9HqrZMbUcyrWXEs6i7NArlE7CZ3icUitPCrPvLI2gT3Gk2EWsmD9VF+b+i2+mm4sF9wZsMSG
kNHJwh2SRGpQH1vnW/TbMrnQK6iMGkcNsCzAk/AEtlg+7q6u6BOcDfubC74BQLN4u6EoGDKpZNq1
XUwmgBACiYdpMYG6OeSzwJa/8jAtvZJwI/5VWS7wF8kQf8lX3+TGOIi7+W+WTGr3N1w8mlm2vPzA
Xsfxooxhe82IslCQg5T10HdekvuIzHIp3puuHHdvl55E38ARXQFpS+zWdHZ0Kwfq+v2QRd4iBeTA
WkWAXqGaezIDHtcgxo93Bh5Y3NAtmRK2f6oK1wihhL2cF+OKU5J2IswEgx7hT14vAsd3vM7fEfEc
JJRhzrDbA8JODWs71ed0HBsGYB2w6z7MJxqLs/SLVU4H9gXLfNciTpiErkVgN23TCvhVvlkHHNJY
86zI5wSXp77yUF7Wa1s3ZkbiBSYYg+WVUCdFUcgwlY+NKLDR3xWmgP9QzTb3sHlckau5YtWUR/tJ
xPsMhY9S7xgXiDM8dFOTCrjxhaDCTRrqnt6f1prD3atpr35L41HgOUy0at5qBX5uluj/LUgLDYfA
InFsdbvPLXg9LK14ORqLcX2FxWMMQt14Kg1Eym2qERuNesnyj/Op/I8EEPRd7mdeRWtqdbfwhAMy
C8xejCb6+5RJp+tXhsM2Dy/Sy8lqph4wi3e0pGRQ+CTgEbul0Rlp92nNhiIQJsvpYZFeivPIcj1A
c3huZneCyOnGFA0IiATejX9opfF6PNNkRB3qNEPABw5ir080yFrFpPo76eC/jrAO+QZAhp4uQ38U
smCDa9gspOdB7xvEzVzr+JgyTpfkkGxTaOwHLCWlGlfqvPO+mAwo9PyNDbVHry4Gx/AreCUhLanJ
/y7zEwPPxbdJgJmlD7U1i/N/nKmO00ABoS7ME+4x91F+OD4tc8RoeaYyenwwCbt8H3PBweUPjDca
/51xnFbS9zUWEh8++c9ID31ij21YjICtDk/NLKvi+vooDRegN5rclHTyTMpnYMg13sIo/7+/zcbB
4gxe5CEFGgPluGZp5J9qxJKhatsoKW3gpglKOSP70nZS39zuMNaPukDGf2opzD216rLWSOfdWxoX
BeP7E3jrZRIpepyv7MmMARWs1PUSayKLmDtff361qatKIaT7jvKKQ3au3IBFVjl4mLRQcYLTv5ph
p071OICE6iVV/YfNsgH3SCwwkzsTA8pzmfdpoz1i+7fqOpgvrhJk3t6+iLCS7fu4x7kaPRt3Ejbw
PSMz5sTBvyKiyhORkOMXES3Xrl7wmOLMaPi43e2X5wccCPpTvA3e5/jmErDRZbgqVsdkDdGC4GVj
/Iuc1mQYOWLXINZW7QLSYX+Utwf1pX/ExMmoZYjJ+9tBFY3NF9pwI30rEE1uG9oAl795N3YDWh/U
/T+QY2RCymTRaJ4P28IkxbDzC4l9EytmJeYaWGaU2y/A4tLzQ/Ap0R12Dza44rinRMrsIWaqkpkD
/Z0W2GksFUiNapqUCBFmV/Iy7lLcobKnDT2O641RG3LGdTIEJCBUyPTulq3PytPl6PWtqoOnWFXU
eUWfLTCGTQNSrN1AnPWZuKh81gXqoNE3MPandAhBE3BdYzrCPlR8gz5f2KPLgusG5wsKAsYXEsRj
SO8ojdqbLtMBdf0pGiF80vFC/5wUCJXWtbDUlI6+FG7QeiknWytejAeVhKripxYbdih24pCwmWk0
GUj5zGzX3fpUv1hbIuLSZKoBVOK780/6V24x64ILhKET+lnoSdkJuhQaL20K33uQO/aMc3hyr9j2
+lYpIYvlRF6DmLTJcuN1ERJFvbMwhHCuq5b5qvQiQ1/OEnsMMdQJFLyYtL2EgsBG0Qz3DWlIrrwO
99gjC1E7iKxcdftrsR/56uMfxPs5A6XdbUImXHcFKzZXqy52weT4hgG1NRx/GuT7kzpgRNa9XMWb
ZavIDFiYQ/ecz0oKDQzmr253Yj2YaGONylnCDB0IL9DYNDjQcmHGVdIut8VcxjZ/aepISf6/yYYr
GJ75jUQNB71mJ92Ny8FOMd4ukQ/Ziw0wTa6dCNhq9ixuJ9wER8+Xx2eh142n6GOKqHQ1D3CVOG2g
sA3qMqj3gDhwixM2KV/7Ma2vPrDyev+enGB5yZhTSf46BJnFtLwC29wI0KZlHc43JGmeMUYaBuAj
B5SjE0y78rXaeLiQZ4ZwiJKcxTs0vpp6NrlxBK0/qrZY7kA3mmOvhTuERHG1FzBxOqODRwegg1V2
Vhdhnd1h1m1sDcglhK5y4BPno/uSSV8NcoiuFLXZ+7vEAjZram2z7EItkw0dL0evR1o61AU18Oqc
JRyklwJt5ZnxY0EnrnjDIJHO2s0YvMbQRPOwSf7swZ+yPhzAA3BEN294E2hwXhWIHg3hiAEao4tp
QZB+7bRXRaqEMNs4Znj+7KoUrpVlTM1+OHHHpLrW274fojqraQJPk3H0aXnbQv/enYQMHq+o7zNd
WdrMCAuKzWEBKk7eoC9OO2Tknh6WrtWdeBpWKkv41rzLenEp4riNw9MNe89XR8WYi07GQXM99PZn
on23uaqfX+/VZEI8b+UK2joZKnfjtrKDng2Gxyvr7H4zjeSCKUcPh0bSjNTg6a8j3ppePnIz0tg0
wSmz+cg4zi7qIDVqcMY5VpWjbUBvmFWw/nHbkBGmaw2beknwtCF3+5Beu5VMYooLLQa2xPtEBJYa
WY9BUtRbNsAvP1O/dEWI6Lckug78hoEBGkZ4/KI4aswtkgMHE9mocjaLyv+oWIuusDTc/DhQdyF8
LiXua/bjT8CV97Cvm1g6YO2mi1V1kCKFq+MKSSUus0e316S25oSL0KbrctiqympsCuJYtaGW/2v/
jLm9w6nf7kSPxC8dgkEEXKNkaYkhCh2Kez+lSx4FgUzm6lpteaI/Y78GulNw5R6nb2tAEh3NnWw1
7HZNm5VWgpdORvrBFHz/oRKqEbjDjKhhzChTgWy8vDg5JW3lxlX/U4PXDjImh9NcXzK4RalYjsED
x7GVkhGDRXmuyUyQMSlXWIJuM90RcSEeEQGc3jr9Ksnk+wmAvHzvLKgL6KOwv6RNge0aep0oZpJH
mTAglnJNrDwvBQpsjb6z1sJ4WwzQjijKfR6hEqfnmpdaSNC0fsw5hU9IJMpYGTMYonCwhhYqyseq
p8yDoLRUgQK094TQUc/Jfe/q4t69U3+J1YQZjaUpsvkNBu6LlydaGmqrh5QixsmjGXS+vtrh4jAI
1UGjtxwyHgzOEURAhSJOzN7uUhsIV4fQYD0tH0DjNCQ0fauoF3PShQ6Yk1/IGARt7IJU7CUNK/uP
qBpe+2zuf75m059G9D5JpTOXNM2smxNuMxKYDQUF7iHAhMtAk6SmHwNVGukackvy63n/oRkpbPtr
a+nmDY1eWjG5H9m9HS5u2thzLRiwNSYVd8WoKeuUZ5v+1xoMAd5imQ08QotvhwBSeUPEiKCde70N
IESkIEcygSKWHhLxiFQtzOVOkgkOUWrYvNLytltHAdQCJ2NrPk4lzjiid13aaFsAI3YfY0CrL6Ih
JmqUEzXdRJnLsbqVog+QSF3f0ekR1Yw2LXdX2MCzH95QlCpctpOO86pgDv+OFXPl0VlgOtGxi6wB
aoynOB1Tdtohwd9bAk00Vn5WL7WeuEyNWWsPNF0K/u2Ym/yhsK+4mwETrxGzgfKgcIKQ1umMNwi0
49XtFSDdBqdZ+p2cBQhiS1aIP+Pa41KyK0BQANXTJk5YbVOGd6E7si/+0/SfY3IMj1yfGw88kAX+
+HkonmBSKGjg7gTRbF69HisD6jMaj0H4mxECc9VDSfrmL6H8vP9927QGp21g/4ABiY22PHlCX1S+
YabcBRE3+5ZobHx0WFWs3Q+Pl/k4tgmT4nZ6rLKl+JbkzKafp1t3UJuXSWp4krVzmKpQYanrUf57
s26W0wxa9p0tC4mU4CrnmKDemyeAdQ3G69BKgPuCZl5n6kjjPW+uyVgheVmy7fq9txgyyRdtPTdL
t8eXX52ZKFbaDkUBBh5+E115NvYrSEE2bsTEJpm6PRfUZLOIqqOAew+42LuIkQlY++VZShpA3WkD
F7vc/LF/FU0KmwsuEpXEPTFpAEIlQrMLt01UYSeYIsXWjbpNLXrfY52XkpoKOGhmKvRWW8dVdbPG
TrtFzv9IQo8JPe2+NeXXiY0VMg730o8fDVcqYBOnHbC1HyanM70+pbSOjab8JM+DpFXE0lgy+QgD
VMVdpntaXKeMv/8J2w9t46TCpJ7sU/y79FMePYukOJ+zg6I5MX9FvwmfJkYRPkwZ6f1/ARkGYtFz
8S1JDK20iTaBMK4dUee1i1dFxp3pcbiwktEf6TO1cEBGFMwejsj0dR6g0689ETGUdrrNWuLf1eQn
9ipou14B/rTAVdZu1ljLBxlVXqFJijppSHWm/LG3xzZyg/HdBlClQzBRFwUJXCOAVL13YPlyG+tc
gf9Z8SWDAIex4Vuzn529xGOxkum702AZxP8fPR5tf2mlu99TTaH2INpHYI+kKY8aAIcvvOnMuZH4
ikHsJKwre/KXvr0n5ay6KmtJDH9lIbhym/uUCAiQsuYS6+Lu1Wlp5j15k6ecA8VkVIOQM47h7SV9
uSotJFDlywbPRXg+FZw5FyHxnh4EJ+tqL1uz/IztVy0iaZMDEVVrETsfLma4FBBHWkaS6sgq7KHT
kEAcN3UW9paicgYA1O6xNMuXywvxh1+pVwH27LvVKOVD6JlyQUziLiT57sVF+Coog3nl7QJSmZwi
srE3bx6Fxeml175hfHKvKzYCdn9g+25G45QXPQMOK0YqWjNIzpCOl5PVeGxCFVlBz/dujKabjkcT
QcdlKuZzcMnSBov2SCc0y709WG1giHhQBGLqlN8357keWV1KrtqhDTMl1tV42dwpmHrBtX1sEbh4
h0AkdkiArfLKQBsj8MBZYrLvSH17Vj5QDyHEJHlYZm1kVHLxidAGMA1TCRfIOoyUy+7QpqG4I4pg
yDupysRjxgBFZD2Ra3SFOhMvKxSJke3hJ4tjeGE+aRkx3a83aDM4UYMqxdZ6YjL5vAPvWGKlDMSk
+IAJRdPTg/eORwN75/OwuChG9WPUzTqfByKIrGN3XFhqC7BEllkSLO4Egr5Zb7goVaUnEEBQjGwO
CD9/JBjTOpDAczwQuLGKVtChhH/GCJCmaGHgh6hbAHRdBcV+wfG3gUzaa04B2gaAc+p+aN2CUGvR
aputl2HxQ9KcaW9Vwt2UWboWct1alrR5U13Qg8DGlEsZzd/nzscjohcC9LP6MqdnfXDaB3Nq3fnB
VFSHIN+SUVDZxvG6E8ukl7CRUO4sh9vl1TKpx+r1DRNfFYPjiNVxABRRK1wJNK77YnbiIEK7FLX+
4OLriKz74/VxFJHf0Xy7wwpAV9jCJ30KHbUvmHtK6OenzFsx8OrofBP8O+YS/ybqgKpmU8JShDkJ
LzSxTnRaZFLrCYxFV8dh5hD3hValZvJotYf1p9lsmojnGKr3HYWo4WaN/1WSd8UzIkpAFesg2AzP
nIV6OEPjsyQzMbqiQSJppxYLgk0pb5BvAqe5SbRZuf8P+Ax7SW3a4FdaI4XENjX1Sd561p0bPlpG
r0s/M+sgMOApjn5FaIrPddiXPfHURE7i+KOf2VUYsAQUPlRFrJejTLohLWsxkiFEClg/FBAju7p8
KvaMH21I811LmWZTDdvsA1hjIp+nmG2ndC3fM8IPoYXvkBHUTZHneLXCnZNIklPJ5C8vhLAkzS96
Sop/0CBfnPD/QoG77z06pNN0evlIAQzeuOA3j7Tq0qTa57uAQFChLFOis91oQCIcS9zYpV0WzW8+
BbpCu42/a64T+Lo35KG5oJtfmYNN+jaDy11GGKymI0qGIDOMeOmAXsBYNVxtjWvBG7HSpnkC4MMg
C5EWRS4LpvDKJevgd/0RzvlOySsRFwzXD6ZMbEngH9nyjj07KZWuEmtvGDdgJFqhZW6MMk2XM6KR
jcVipnBIcxuErl748fNmePHxJFZy1Fs9CUVBtFX9SNm7OyB0310BN2oqmOqlR9k6m8ASDT0HoLMf
rqq+sqz+q2QlchvxsxdxisqQhxRdrjmpYh8iwrMbZrwNS/B5GX4TjS027bbhWS0tkSOjjPyBQWmm
Far/Tt48tjIWif+L21yYUIUVZv3QK8xhynbvUGtArfAIcctSHoUSyd4XnE0aua8kFMSuZT6aL7M5
2m1AkvYcq5aQlLZfSBcrqRjOT/97KDrHBgx2u6VX1o5LYwvv+qDcAnyT48HsGAZBeO8hG5JFccpg
L1P4J4wkrQ7/7dB1FS7GwYn6goZJuQ4DUPdFdAj6tb6L/Lpro+4tkyNDTFStBSsFIV5GvzR9sv5/
odrwSh+gqywu5p8CT0Az9mcIX/K8cibwVzBnb1r93BW0oV//2HVeaLCbDwYn4eBggPfHLm+6eBby
W9q+oQ4e4FjVnyeTUhUvwu7fcJqzajycKUIq3p/bQx+DuydF3q/zlxRTR8tm2gX3obolE05XCzbP
0I3cHHUgrFqty5ZGi4f1uHWNOvxFV36keBSM3THzdbYSb5GlHMODkGVcNZQDdIBkQJSErLXz7Jfo
4pvMbuEZ4jpLXaiLNWFzICYcgYhDQOCQbyriFk0ZHNxntcLbMXKjHPaY5gC/B+3su+wqINKklD+m
CZ3L9cW7v7hajO5S7aizogFtUVkHSn15X7Te1BdcocFBESbn4kFoNExQ/V0DwMvUGiAZxgmMyUGb
DrDwO/9DWHKu9Ax03LpVxtx2F2+Q0Jq0ZR6xSj2rHPGxUxT1iLxqObtZpoTUBDRm3Io6HmgAxaWN
hzqowcXgZ6o99KDEQ9a/oStopifeJzBTJevZp562qinN0fJvERsvo0vBvdMEDv1sWOjFnL6WOYK/
EOfKclc+aliSWTXzM+uxfn/K1nUd+h4dze8WB4AMaTO47dLIE+dpCHN8ON2VDUnLHZwzAfPsC8j3
zfuhYWF11bwjwK9pKyYQXn7+Rzp+C4QsF6NSX3oOXeUclzRpLPjh+pyAnsrNmlBPBjhFHtOFYj5K
EVlpACddiXrDklH7HhrHjfJfWkrX0cOWfTK2KrgyE6dZydgVdd060Xw2e7tTUPK7kzkLhEJNn6lc
r4r9eLeWfGtKuvahdvDqlPRsAiPDMYSmx7iiwTaDk/ZM3cBmTDG/F6a+UjIFTmO2fy13BY9DlFNR
w+zg9/QUbLn1UBDrdAva1A4nuBhQyr1vuHkYYI1olhCQkgT37lvnBvo2lzeaA/sPDWYKA8HvgAcb
mC5Hv9At0CNZR67LKmpYNuU/K2epZAmYDJb1X5l8koQPh8DXZo/7FE2//LOOuGrTbWMgAVmN9ONN
KB/GylOit9R7qtQYJgeqgOjiNsTSYhM3mOJVUIZrCN5k6SCH0UdiPsfHQWuJZgKZMx1eZ+trxCow
bPLWeBeBBoe8CeJlPhw9YNHaSRYT3zHMuPDaqeJYH85ZgMbjB8mHCSR1t1z9mu7WQe7dTw5lMVZX
AjY0uzFjZ+YYlOkYx/6JgfbEAUdX6YnttFmCQMEBCthkV647y7SR8MHW+s13QwFBYJn/VmEVaOJ5
nPOjhP/WwQBCPRNmiL0iidrlEFiWYX9W2qamFGglhXcDGwtC0LK4ij/hlxvZPrHcDdTTKqDGR5zy
xR7T0MBA+IB2/rsS6XBJtpJjXrfXRpgR5kLNbHqFNT88t15z+ZIGy+/R7RTXsTQqUHe+Jcm7SeGz
64MZUR9CNfqNdZHaihSArZQbPzJTR3oh/WMvGs4/F5B9JMSHkL+RmArhuaRG1UozCX9SpXE1YaLX
ji+IaARtONaa9mKF308hQ65whbqDOXZxcdh/26olpkOvgd4gG3WMrMd/5jGrjaGg+LCaySfFEyM2
HyBheUYE/wASPpDc7sdZIweyZ5sHz8SBmgdoIjF7+nrFS8oO9IJ9RDJzwP+AfaFcy5JSzEzxA8xO
epF1MIasteQz1FUzfQgliW767x4gybbA0UOqihPbRmaBy2NPonn3j7VWcZP+GW1dPN+6fHGzH1KF
rQSsE00GJby4R/h2OI4YutlPEFRH6BVj/KFPYWkFN7orP+xiIU1dCQxbLYhHAeT7bjp1nMptI1gf
7wzgIOdUgw25hptTvCRAz1Op7kSup01ErVqtsgnwo5BeObzeMxCco0oSN3dx+ErdkRZGH1SZZ3nG
YsiQvLu6+l+7qVCzmlUF+7p6nwJ9405UMDCGG1pcNFwq8vdieUOMsvon7n5GdnYS0LMsHkINV5L+
pwEWyffwjMIizFeAakIBQt/rk20SrT/mQNTZoO9d2hexrkNvoFCdLjEh2fE+iP34myh0VkjXNV+j
gspFBv8rwuKmLtIbRG31eqT7mRNV+1nFDpm31BtoH5nE0iKE9uA6I+pr0A6QKfZPwE+Wg8po/1BA
LS81TyrevTd9u81KbDhu4xpyTpC0bk34lzed2LoxKQe/qSLE+b4rv4Y6DvgoZWRcGl2wE5eCBKGA
yZcZcSId7fbI01XbcqWWCjGk2ggjcvD++5Ufxn4UbTMDoqkUjZkzG3NEplUwgWU7NisScLVLMRbj
nbIX8PE0pSqlthBHNSrO05w0z1YPs1PNs5MyBx8h+AESkT0+73xZ8rYLT1Npy/uM6NjEEU1/CL3c
S5nMR+De6n5pc/qtXa4yuDT+Ala0au1LV3teWAl6OEs0MUBSAV5ZSkuHTOuNGoP1lLHhw55dDX/k
sPoaYBx3EvAueH9RqXzPIMT0z7I5adsBc6lwWZ9cw6V9bA10oP7z4g7zlegJZ5AJInMpBv+9gWZ5
JcciB7JS2NDwuMZ0Y6aycpLexISQ50RvA3hCJQvfdQBmwXpwAVGrs7uo9vElZOLwZ/2LigdchXyE
URFitb9gm9ROkvXPeadrJ6DT/6nBu7eULxS7kNAm4e8VmyB66KvbmCcbE3S954gHEmDraoyup1D4
ClGeQrfqrq/SxhQb6WY9OFjHBVkbl8c4BUGhYaqxMKPicqqcu/fq2o5VAAv6KudIqAnWe4AOiVIC
G3BTLhazd+6xh/a7zHvrOTQ3E75WoYhBk6vQ4sjKerjhXVYuaytkgDpOu55xfmjX/+LTA/MEiTjA
/w6QSR3DC3oljV+RXS4GcQQUdNJxkF17D37ZzVV6qe6l+i07Viymnu/9x/I7Fm1Ttzy+WyLK1mhz
icOvUa9KNqsi4vKyKNHEfnn6d/X7eIwumvpBRlWBYljrVBQeqMjd4FFpxhjA10SzmIt6z2F9Fg/Q
MQ0F43lBU61uY2AfnxAn8XiQ7jxHRfrsO/4VKq76TI2pE8Thq6m8NAsXv5o4ARLNkkeLeuH/uyrT
8x6+kAMHyDZu9EylCRoeSYhuzkift5t52QLm3GkOlfiaerX78EaYBN+PjAlezs5Mi4ORIhyRNNPt
pHHKBJiidz5Vy4YQMCAb9569sPSLbdK/HYrWB0qVLJmXwEznyBFvlI8cTjaySm4mWhDFpkUnNp5s
fZZpgyaVz/9TGjEGUeNgR4dB7DYd0GD7pBur0vZpmJUo8khH/gIht2C94dlhChR89HAbG5nwMF8V
/zNO+3lkgzVAGLA98Nol+pIp+2wHQEXb+hStFDvZdSVpwX2BM2KkKZci2N9DRtLYRm0ukWZLLqPd
M1q3LgZ+A/pQPPrVaIACcv51bJBAH1RNqjGK+aTc6IrpfdCyXNGvhRBB+4NqFraAutXM5PN213Ua
75YEm3Gt9tz4aqcx8doUt+zZU/+VK4f71ikREW+TLo0uhtHvMLbmkeI/G7588bbrksZ1cLnoV3ip
gGsxo2JGfdb+1U4q5xWyQc8iTpok1WGQ0lkvGJDFrSvc5uxGlFebDF52Q7Q0pK/0vJnX2UHR1FXu
+f7dEVcT9ShOcf0YlM+xf9J4zWeBBoyZn8b67zs8JwdkCo4jesNnpMdCwq4Zb2T4vt/r8g0Z2dtj
j/fYWaNF/pyoFTCzTSx1s0PZV/qbpEWhDqoanoTwYo3jX5kWsAD1HlMUgg/pXvNGZGev5OKpL2wC
od4rfrukKBB45RjpjCyYYGIu3SvuP0nSHifMPVRHmUIboQbrScFkxhMNk3PwGY4G7Z9VfuRvmZA6
+DUkiyEYwJ1qVo+Vr9VEpaE+e/LRXo7pfx7Y2qHDa14ztEA1rq+D7tOre8fsp6ItZkghRxzrIv1U
nR/ccw1fcTqvgUQC6UJ2L0QgYXRCjPjJE5DWUZMEEfuabl+uBYOU3pO7aPL7tymjmkCAA18FLB8f
gtt01Fe43xHlV3wgW6+/dy/54JHbZtGvPhdkwrFDtBjW8oCE5m1FZqmwu18Z6Lb4eX+C3HmVs7+z
VEeM896Pv/+ZSD7bOIC8J3YEs8NO0J+Nrei+5GAPjXhxWA+IsVbJTQxyJ7J0DbTsNmV6k5hLORPP
ZpBXT/1HHAMmDH50mHtX9udRzAjHSZhik3/G/5KDyAoJTBCV6JoHxTgrIJCLWLF+JBPeVhmgsVle
ervEqanUuwjoE0H9oS5S+95uJx2cxswBpkAYH8or80hkSoXcWSdrB0LjZpnbEM64TedbPpqk9sfd
gPEAcCtCuVM426UFSAGrHtzCpmha5p6Qxv+8EP7KEZ2R1eU9OcQ7ZgicBAj4tgxb7oYIO+AByOi4
Cdr4X3KvtBgz5+A94wqmXwrI23ZwcH8Cxu/BwbRyb4ZXqPnd4tRvTo0m8O1+ftBW92kYliBYEsEq
nFpJ37ZNhpQsPOhz3O29jtJEcOuGwf+uM0LzJXYwh7wZND5VxFrt06lfVX1x9A9KE0wlkMIed/zI
pmPJrdcT2u3352hQa5x5YpC+1aUgZiFFSnaAXst2M5xiDPtNtLyQbz9DcgkYHS8ftR/lxgJGz3Wp
nBP3ZydHNAPWZ9gxagdETO3nccdLTuWMMhYmgFPwx4zeHhzYDq3fozNOTsCNhyZyBMBI8Z3xd8gk
ag86sTNDUEFdQVIo8hbadioe0ZeyQOB58CWp+O9g9zZmB0bXpV1kDGqghXHb5C2k3mJFvp2jzKnE
SBRUdSGTZBcRJ76nWH/JfIxkGo7f/4CyKLiWh7wfICzzm8p4jDEvZYwHniR3omadRvR1FBBJTpKF
L9IYtztXC9mhIs+3IHDaJv+uYB7oUp2DnaeTCxfsAoigGJzLQ2SDj6ed0FjKyqqulF8XX47KGjzA
jqzqB4oYZNIWFJe6nJLvNuE/ESNQHZ37rdH+3hgrmitC6+24TG0j4GW2swWpcJA95UtKtZ3rq+Cd
FCcVDchzi9Zn0V8q16MYmwszG85Pzit7+0hyWEEXE/r2bh40lSL2BpgM2HzXK2D0pgxCNVZZoxys
HQ52YcBW9wSUK3I5pM4F0OW9ZkG1IeEMgz6vyomUDufm2l5xQDKjfYK/vchPw15s5aboXEH3Etqn
0rDaoYMJeApmAfQhuGN2oH0oBde6IWhynTNfyQ0O4xv/EE5rO3thOtDT7dqq3hrriX8K/o3ZXuBP
iPKVVLemNGqzZzfJ99YhiMAe/XS5gZWNjvg9nNouCEAkPHg23IhNjvJe7WihTxWqfJWShZVnFACS
+DbaosG9pQcngdvZ6cH9FKjE+1NhZZwRbjshERHErKriiPKxMwRZycEcJpdB7ikFbPOfkQvLnSUD
dUgYdnd1CGaJmAIppvNcJvPQYq1pV5huDQfwSDHPHIG6yQ4Yv5ysK+G1snXzr8R+jPmXbQP+us8t
wP7jhK6LM+V2smv8LRewOh++OgWYjZYr5qgrqVjYQL1ams269X3Bx/eafqzXLCwwRyz+s4ChQYCT
vcfg4PAsSYS4VW57W8c5GyDBqPlzIH5cvrnAGTbWMF87gOQHOzicw4M4ImnycbK0A4cq6AcjtBoi
Og4TsxZzdCLlu+iNLC1T/ErSTMjGI71yCe9E/KzE6VE=
`protect end_protected

