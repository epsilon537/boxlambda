`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fIrCZrLebFpeq6OHp71l17OSDRkEgfyaH6BXlsXkYKgIB2q3+YIRxqsdCIM798CmIG8oPOk5/rmn
xFrPf6TnCjG98pQ2McXt6REwykUy/L1gYI3hJA4bHa4nLo/m10GwSd7BFi9Nfw+FjD9pgb/A7nHZ
OHRBc4fnOqeR4fw+QszisMBbyEvIqaCs0X8PEZPoaxnDFD8PVGrmPElBfovoeq+QBbXhIE3FmGQH
rWzaIo6/3MmFBj+cUORwNfLFmjmZLhTuAzpJWHbWeWjMO6V5OZLFCHTA59WnIt0EEAJzdmkdPDdr
q9pjbnJGmBgORDYqpsgFzrmc5WPcu1wJMLFWgg==
`protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`protect key_block
rf0bfkEMrERhY3gybybh6vKlkfa5na2DJ9i5+Efxmv/IkLTQ+1Cc3GktrybUt94IEBwCGV+EVmbs
OFw6+8Oo0zsFZ2/s58XJKBH8CMWUkutC97pM0SrztIkcG9fxB72WX4paQPKIXdtUin1gDMNCEfE6
8HBQhPrIugfGSJZJmAHnJFan8jiClfrqkEC4DazKJeT19pTJfrFAkW2BrBRGUN/BmTuqjQuQQZlq
+K03rhlvb6cSup6DiS6x8oew8pZsSpUawW7+UV4YKB3QssMFJhsFnrYW70oJEbgdfc1CL2FuHpSq
EXhMDjFM8lsY0/q4llZeN2sI6Ne2S+j2SWBMRwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fWwY+O31wo8boyWoMujkvtlEQ8oErLyPyPELRqCa8sRyr1ZJguYo7I81HS68sqOITUVKTWT5sjei
6aEfIi3rNg==
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RFCpBbphraMJUr460M9giDgmUBblOeMIuVgtfgSPUEL9aBVXY1sMvIb16fQkr1gWSRV7I89ZUb3h
dCjXxq01VpyYs5TVrVgu4Rt3s1jJ9SLBAB8KMyp7du4KYUy9lX9gF/pSd1pvItR43w6MDaMqGklv
aEOBsYRQlo0hbu5xCI/LlKdZdyAl8IgcU0bUTmuFSItNLq0v3BET+hOBKOUzxSR5enYFOZBgxy9U
4z4vQjUdgeoYNRZuxrzW7i87n5vTjiAgkC1BUeXbRlpFEQPFFy0n0VKKYBqdSTv16+6U2J0lLPTs
1MjZk5RFnrfXxS0MptrIfJjEDJfpme2NREufhg==
`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LjjMSTdGKUXjDB7Btixr3Ysx5w2vJ3ck+cdm6w+zyNO5HIWDBFLJw+rRwxPbDGFGcxJ1OG718ZLZ
FYuWesUeX09ZuU8hj5fIOk/VIWV2LRdtZSvO6kkimP9chB0p10IKEpkcmTE4Hrli7lFAMKkFneMp
tri5yQqjhE7pwlzEJnLS49gHIzvpdKH4ziHm4HEkDVwreI2/Enjm78h+kHudk+HoRLLw0EmUbf06
GUrqKO3QTW+8kfbe1q9jYX7uJSPhhIahnuIjszoXfL0MfTLT+pSdw/iD2XX8FqsO72v2+FRzjDvV
CquJDbdElNE4gnrSetVZDN2p89vgSlvlr/MbEQ==
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qdkfDAm/sV0V+ps2LNv8i93DWw2i5G/PhlErK+HTD68kNwnVmNopsqCRVchV4xmzob508XpnoDwo
+DBdl5Gc3K3fJp5vFgtWVDT+filTNRyEz1bv4gIcc9SKje51zpMfbV180vfAWFZmpvnIhNLjq4vm
kytdkRsArwN0b/+6qHk=
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AGaFniwhlaoS446lmm6jbjsDCmEjp9DcFzWNJQQRv6opm4fud4JgI/jaX9zPYnTK47nxSB12doFl
FvwKpl/p4YIjfWawxQZCXM1ppKmsn9t6JntDgqPk6xxEzIYRes4BorMxdrppID5Kzl6xIhPH/hEV
7aSp+DWW/1pwpkCi/WXIzOJ3y+/cOJwoOYlg6aWtYkKXgj1fpCmPNe1ATlALR56iDnnWGekJyafD
ZRY6V/Upn5I1uatFEol2BGlIYF0Gb2rLthVQmjCbx8jvoic9jjmEglsOM633SNzsHsWYLgtJ8xPx
mFel4lECx11ddzdUCXhSfmyNB4Phh89QjjBDTw==
`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZjtFNv9F7MZ3G36ssAmNEAlWVeJKGoZgq4pXtkfdLYfb6lnqOU5IATzw5ylkTlUdny2I9WgmLKHg
gjL4ztnnMwdXtaz6o6FxRierJwdS2JAVbOwy5uMzEEvCqJMTHorGZ1vBqAGe/K40QM5jmbK/IKJY
GBII/zbHy+U0Y18iYCBXrltQlzb0SRN6w3BfYfuYhrOSPo3IWwHzOOlfOME4rhg5UhM4Lh3XQU3d
gQ8ZCHdfgb1U62ryrlgfVawlI8RPYgG7CsGvfZA4sNQNKOmun/34lDPqqubwsFM0UupPigMyzQFD
kU/oShz/PYxb7Zg1KRdIoLIs+qSMOuyUXsAoPg==
`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cP8gJK9xzxAYzyae9IXC73m0/r2PyMa9/QzasBK+zuezTQYT4pjaJC0LCyhaIDLLULkiFw5P69Il
qX3vx8qgz7UchElP2s8CEwtRwk7hcS++t1gQjSNFQ13t6Oyl9msTdyfoPVazHVDekuyVE090GLlg
/jdpIq17WNJ1M91vhGY=
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kHKdWYyTkb0MABsxTO+l6zE4mFxQWTqDTKvtYpqLCmp0gtH+vBrpXV9cUg5khg2BTSClbo4s5RsP
CmsVWKQTFsnMpHZnwkNqhLnd//cjZCP5xq+NGdUjIVN0qGJc31mj4tEkTYg/Kwe8pyqYA41YceV/
rC1TA93Ur7Oc00t1nBYTsm+XE+ZeX1pAW7HjfnrqKbGiXjjukuTgjYvEl2m17JdSMfSBGg0pK15J
sVy1q3QsAS3mb0m3IP4obISoFBN6GYLcR/Il5go5DnRF0Y6X32yrBMynV4HVULHQkfbzZc4uNM2d
tLClYwAX4Se4hL2NGVsECgNm13Ueqh+iDzBa1A==
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 53760)
`protect data_block
XKDV5Y3Lt613kY738mjVQx9Sa4kQZUKquJQxsOZh3YlEaICE238/EalXqQ6g5FjYdahx3AC4tfhq
olGxJMUoSQGQUvD2U/84Var6I0k5nm/dasWSl7fkhGHp7bx8Dted2nC3wCiunurVBNSg2FTx5ndt
cVTXHMJHMcZ57amD3As8jWlO4Lyb0x0JhastDoWJm8otKxPDNcvyNyYAu2Lv/cJ3tKyilmnQFp/g
O4DqwHQnwpxLktpS0ja3IlSZ8Xe2AgNbtOPkayZK3KSLQQo2JJxtOLU3hPe/2n2l+eXto1KUn3D0
4E5F42a2LwdFKXoCxNOlVxotk0AKucS25eAeo9xUKl0P4DpS8XqdcqT+aFzaVOWB/sleByxYKSKV
9V+KuKhd6sjAcXTSacuQSYyW3IsQTVql8ZLu+uCBhEIw7OWnSX5dzHSFFdCNs6WaM+jrydwvY9HA
8lI1q5dFaP6zKEYYQVtGD0wna0B+/apR8lyfCRaMBrr1OXOcy0nvJ2PdGCUKVKJhDBU2x5eoOa3h
dUKkTPetPi19r9QVZR88VpohGQDT/vna1P/Di8oq/w3K82b8xl5PWMIGibV8pqOUpGlPYQ2nfWvt
OkTIp0+0UBPKGszOvOYfve6qAOn6LSKj0wGypFuPdKfVMT2ux72mpdqO2gBRrvCuvdkkkTD8gdav
/J0qs+Ls86Z4LdXBavufjZxkoqfGjMyhI7Y07rfzbM+BQ4c2hqMNfqyCi2TnyT4KcJ01FDA8hBYG
GLaxVytAXASVC2VBA6ekLwLEGU+ZiwChxKpGcXTAptE/7Doq5zz2miL9B4XpqJicsGl3Bdxr2ONd
jPRQZv3moSG7q0b6VZwcI3IoS/bynw7QSVec6oSsoA3DKWxtdXT5j9/iU2w2SxxvvDCt0ZY3xEC5
NhzcI9t71wT/RVplZc76/gZ0qTslTWUEuDIKaGKrxONE5pLQAMCDBLNapsTmvIqSijbF15G3pH9z
Vy733vb6LrU3CQT6hVmupVFgt4AqElSjIVE9jGA7/+8wpC3G3npbOIvBhF+lI6RbbYCTGYW/Q71A
7ZEQjPlGb5WrTgFCfOwjd6No8tRh2B3r/QyYsWiJrbNzLUoPJNuDhp6dN+2uACPTWv+VqRoKwc5y
Cmfd5miF6ATDwdDdj/32QOTp+i9VHKu9VB5srT5L/sv6lRCfmrkwDq/+HLTk8yDtdcZRLPBx8Tyo
28NDtfeHFR6nIAhzo6pqgHRphvpszyHOOCsbeHlpL2to2oAgaXYZROOsRFLuiW7DzNuFs9qsI04k
W8IEQZrsYSzEpJBnWNXJz7+wsSINdJIpXJfu8uh+wg14wXHtdmLJq0OhPbpnNpS3VRgmB07/LD8w
Dr5WB9s/VytMOmoGVuCXq6csKcBolVk2q9IushcoQCZYphSg9vhZs2ovwJE8zfetADQ777mrJEC7
uybaZXZ7jsgKHG4719iaUMYkbD7V7HoyWt9/+Oqo4PAzy0FVXh2JWF8ZfrVRk2aV77Jyt+Vu+vh8
dzbuiPxFRjCeBHnqWB09qK7rzMKtUe0j/LubrvckiIFi/cHKxj/M9x/TgQyWXdcYiBKw4ABmRIUc
Y0ljpMGn8QCR1erYyLRZdRQacrRdDbTNhnp9GkemOsRecH4k2WLFLDyiirkgPqeK+fA3EYL5GyyT
2MOGh4H3H52xU52S5dypwmPC+5jg28zFN+KElnhABNH4vdkWCzhM3SeU7h9lw2RcZhNvMA9BDIUy
JS3AKEEShSzZwH/DtwvD4Rz1FkU9BPjUEatEs00POtn/WVnyUe1M0BxTfjALYsbT1PEm6ugxMxg/
g3XnNjYe2xEHM5g+2U79R71kxzE0ctiXKSeHJ/9KyGQjCG1GKgjrfUH6QhaHqrNd9fy8x8pgXmsH
WNQFhVtNTyu99DdjLlrbtXvfucMRrwDPHWznTFnpWWVLeAYlKwr9dFiSronsREhgxP0+yDgLmOoj
5oiKb1sHzNUUqYoGzXunhe6jNYYxx5UJ11CnEoJZcab8J2pWkhZGcxHL2dvaovw9NxZEW1vDCe0v
JYyJ9ibbzA+HH+ppOzQXiLU/hg+HuiYIDmbiU/3Z+v6mKBCml85E07fpdhgAiEbA+F/3DEABtqZD
/m5aI4vrK/gACZqSmE3yDvAa8wdYviV3SsHPFoRcjdhktJ+espEnyf/jTvpbYE6xdYz+Nwlcn0MF
FIrHVpTbjxgRaRJK/vTZI88+extPBPYIv6cuws/QAHIExsj3MhYpA3xhsL+wiVG6HFVVi67viqhv
TzNyGAjT9uKeCr2VremtUlpZnLcO4RClpDUPFQjZ8qoGV/3dhDAjNEWLfsakCI9yfTplciYjvwII
ZNrfAO2Mxbd+s3ZmTk0P00OzqFF+ykqrfh9zAaDdXdw3AzPxT7N0S0BkJk4ZCMCwg71IZboLw3kF
cRnkX3FS4QbRXx0AZavTXsZy29SQ+1msmW/CRA72CCGVzazAcstHsnsQGpmD2tp7IJ4u6uYZfV6v
+20FBSfXQLAr7R+xIOw8E9tP++2jwy82hU7kgmAJyPwWMpVsb6oDvmmb1H+WdO/M3q3XvOhwxMbd
0i4ioxvrpepWyU+264x9Ow2yZ4gd1NmFHSj5KoXWlvGXoX0eMS1SjFM45NHGPUU28agNiZfqzj1C
Ad6Xa4Yso6xwYNertP7tkF9vTYd8CpmcnyV/pUQuI1J3vEGv70Be2AlCIPxZc9BovIBbDAqti461
GDCqNowR8nkHNM131GJGe4bYp2VWKZ246uoze3TjfOQ/4MP7ZasHZhMOFZBMbydC92GmDVmlkZlK
sG35dp+NNphs5nc61//Qex3onFTdVrl+gx1Lr/k1dm3RrwPDigfl8l7zygtEeKHjjEIL90TbMZ0v
AGAqhqPoJvKipGAjsPVcT6jwgnIjNw8xMnpf1WitRqDmfNtv9+0AUki2CvfzWR5YYZTw4TY5MzZl
+JIqD5xFCqlXD5iQAS/qv5/IxmptkMMEpq7mnR4tBdRM5+dsv/oaN8wU+dWGUwolN7i0QRK375Wg
G9wt80v4l8BF62BQhc8HBEIqV9nqfXbJOdUAck8k54foJZtk3bzC/48u6g2OZjrxOaBwnLCk0E9g
KDUjCrTr+GSUfgcY3g4LHJGCUwjdf3+PXuGfluwPP8nBiZc2jaz0DoYvwlK04ijLwwdrLc0T5QAS
otVqFJ98X8XSINEmG13PvTKGDF1MMzkd+62udIhyCWeH7UlKhw0K36PtDVVt6oNyxj2hORU4NLFP
UJMGc9WeU7Nn5C5nEBrMu5KCXy1j8lAccb4uEbtPBA0knffpMnHYzReBoVMX1SPncfGB+6lJKYdT
q+GSMMgEjas2gF1wTMWuoCExH697XP5efryBM/+a0f3DNJ7W/p+SG4HkPftmC1hshS//1xEqlRp1
uLJNiUI9sra051QquX6ioSJoExsM4/2F3N2ndk2Cb+GTJRla6cfKs/agM24u6GNWLUJiY7tcwmkf
VbDpvtxlWW2F6dWGu6xwng7uuS8GmJB1qaL/3hH+QWDljSXHQAX1JSSfWcL3L+0nE0sNzUWeLB4s
RHHavduCCwUt/rvjfbP5vMTk39KVhiPHk7kDcRYkYdHjIdrqtIe1FfehcTAGha6Mys8/xSYpwbv7
KqUJE8qbFwmrf9Pz5zcyNr/xPxfnq4LytdMDa60NR1OxIZCvJckdc/nKhbLJhe4zOyxF4oFIrtyL
kFeVq2+adaEYV6l9NxNscNp7e/EDTD5I58ZmHqK78UgJ2ODloqdCmfPZO2p8mdSh+gp3i2gwdOos
88K86bc/XB+nSMCpZHaIhAM2VXFGtKM9m1uxB1RJ5KWYBS5SJ27iypws17lUEk7cxY1WpB7G+6YJ
k/eHtXZlFWtBYHUTNrkryTbM9G5xLLyZwc/mts1WLWCHcpqR3YmadvelYrofRjbViha/ik7jZGZs
4R0ZIPwhwIsd4UIq01SsWa8YquTq5Tl6Sv2W6WJFFCOfyBbENC0gdfZCeiPzw1wvNsYyfZeB07PE
bHZ5Z5O7Mj7wYM44CSbL7NZXumTS+Ee1buO7JES2Hnj91NWdgKBq/5y7EiaJVzMz4iidcKOHR0TR
vLzBW2gdxSpYe4W6/jURKtU5jaZMoliV06C6zEdzQCZeL3ZRjvd0fZKWebVqv+zMzKZ+uqwU7xDH
A4fMSkPZNOkKZ4dVv0+yDwu/1x6vbXAB2dR/xTdRaspxZkXrWM7KhgcG8LBTlh1gnNOvIYP3Ptht
m6VHFWTX2/yU/S9tfEPZala0nHWO9cqnrtUxchbsIvbuAwbREcK3M/ahBKRYlZUY6LmEhO8wAUCQ
reIr6m7lzd0p0zbQxp/1OeP7RE1rWA5qXpN//SxypoDlyUYfDDoAn+U71kToIBqmjqBIi6MhtTaJ
Sai4DdmILXgBgz3XJzFjm1d0ArCj2qAfNrQJVuOSSyGpXD0m3rwtwaZqkk2OK65SpTkhQRWeKngs
bGoYpQmGkgRVdGUrLBYP9hld8jYIUlSAM2hp8pZSQjMZipNtSssy/BLc3Pnfjav3rDVhUh9g1qt8
/5Y+Qd88/0ONssXlZKHToklr0uwvnNwJLm/KZMIB8wesXYHIxDnJ4ohQD4Ke4tDzNGlJNjrFqzGi
MdnZqgXDgMb/5dK5B5Klyf7h83nopFAOsWDdVmBic+abeDsZKCK5YhNO0EUYJQo4rDxE+iFH2GBX
mdnYNjaoJp4EaGZRYA0fEvMy33D4JjjdL0esIRHo8pPRSz0pGYQWxjcywQf+DJ5IdmELk0wSGjYL
q0Be2znJt+DB6C4kaIIZabjzB1adQghXtfAhe7j7Ku3Z4rvGRpxlV/oA03ipZ0ExGNmeJyNQUZP8
4/txyLKfw1SoA00eH0b0VSX1AeqIEPF0IoKqvrUNyrVlbocUYZAz68fvhpExk9XK1kjVjlaYHo/3
zhXKi2VUVIRPBWZC3uFJkrcim01qbWD7p4rqVBRLs0vu6i2SJfR9t5EMHc7mY8ggBxlQsvzpjCZA
vYT/6l9cXkDAzjvAkXP2qz/EqMtNoYTovszjh9m7MCVcdJdqsZlHLAF+FsI6II/ssThZKcEXBDGh
L7oRVH/+VjtCQ8qDRUS1wjqjzjsp0Vg91GHv4pM2VyWAwkJ+rkcXU6b2F37P6pCqqo4uEIS0VRxq
4x8eR/agnlpVeaphGAhAF6+Q5Wz7cuOQ08VQex1MqpRiKitsw35vhNBYUY/pkFPVAfiCxkgi1Xnr
zajZsr7AOSzm3L6YigY5AwlUajUcyGM+67vA2MjLjABK8mLiOK0W9F2Kh4Xtybi32tqBTvK41GrI
bxXukHRP1PDAygAqhvNIFivoff1LWtKXmTI9BpTRrDzqwDkp0gPdtQJdY6FGJVqv5JXEzToKPNaV
raypANZ56N7SRiykXllbGy5bnYxrFXrRaraa9EDLjWfc0ya6uAGulZzOCqnthOWVjannT/37I+5y
MhXHOdqq1DREDM/qY1pHrK4EIAwObIucP/QFgZ0gl0aMMiCTWEIUpzPX/FkvBCwCDQg6xqSxH0XG
6+ju59438TlJnMOtDi8TwiAUBSufe/h6AoyZqrYxfvChUN+58YzQN2aKnjeyrM2AjkCbEQB/Ogj+
WD+9b1RBUQ4Zpc0dAdqTBephjnLVzsfGXNpHQHy6RDWfyYOZiOJuHfBxWmaVEU2NF+VY96IvpEa1
O07Ys6ui/CZkAGZpMiEj+TvMemS+++wrPokpHnvryBAiMt3W1IWMJGllCihauqe1n29GavGe29cJ
EMtNDjbZMxwHAmg3wqzElPW865JfL08kVkCM174A03IzHB1oh+qvYlHtZCIO8yKc9Uke99DXhCW/
6yHBjycW6zoFszgBTKNmLrdtQWc1ligibtbuZ0amexHg9t7pJdOiuM5ESznYKanQJdK4Ac75MC8V
306P8zcb0HlQc8gRBUIV47dflh9p4jlG/dN0VXxHH9zr6zLlyDvi3hmaaaMM5LLH0VdHeFM62TJX
eqZQ80ksZhbQla8D5GTePdCnmHVirGf9U0NbPh88Q7l6KlVN+jNu14QbhVrIFVNuneB6FHkPtmCa
97HJTRLQoP72Pchfz92EBv0vCftQY2kJ8b8ANQmjuRZCR2ZszsZ9ldDw3auG+mLiw5jU/bu04rHp
KOcX6htmVgTBDTheYDmx2fSbMv60TA/Cbf2WE6qLrzTtnMaTGaFvLhrzqPBXCOIXKswObCscDIyc
NMwMj/SOLN1GRgbKpg5hpbz8zvZoNoaDrxnakRML2HuPTplgtUG5/uqDS/uAoRHKJ30QfzC4dMN+
60MDAkHDNed+UCFmdZoH0KdIJ+jYv8j2ibAmTFi0TQe/NFqBKCijhDgue2mntIZMBz9QTwdtuTMl
5NK8GEo6IAagVzNveA1wXHa9YNTWG9n7x2GDrLbOqa+jShOODZt17MmsyJiWLTUuuThf8UwHJJ6y
Z8gxV5MYfjL15cqAJz3rzmBu3v/m6L57a+gCLAwzg17Bb1c0TEpvhSrFucoWa5DtXmLQCmwzeZsp
wOjJNjLG9upoQtiU1x8nHfEcBKWchEBvpA9iJ81NoknYeMELhhHxG/bM9MguXL5594kooUbSRGed
Is4l6Y9rjt5fdDh9jRD+x9kqxEW4wMJPTSA+FoFFpWetm9oRFN7tdiTqTl20kN2YYY/nLpXmTmnW
Rz6PG4dOY29U6MWcYRq7TfyAdVQZF8GFkk+JCEXrzzUwbiqyyoygrh6avX18bYBSomX4re6Q/EaJ
PQossWipYdsZQWbRNiod3Fuen7ukG/pFvASYUE5JbXGurULIfgIXUQJiR/HGeFKOk/SIxQZ4dzJB
RBWxtpq0NMfULOnaQR2RNHef/MS0n8DHyAQnQ2Mic3iJGJ0P5PDesDh36rQZS9fFniWYW5FDX8zu
PG+D0VB4vF8uE8jyA17lA9rDpRAU06gehldaHAJMTVCyCU8PfzMYqiM3VuTB/XPVYE6tKr2d+VrI
B69rpo3TuXyWhDCItlf3b2rciVSM2odei2i1GxrGkQVOYVjCAe3ulQeG9f9SzyGrF8DepAxsKB93
qpwuh3YLWDB+1uZeCwiOW4ukzPv8J6AgONmLW33ClKpeJbi3CPam03ac1jyMQ9X1SAMVFgbwdpp2
tJ4i/PJC4FRNBeJAzcxqBLkI4+WZ20Xk4DAF84c/LLHilYeW4hs/MEHK6qfhj74VcSuU2958cx+Q
kdhocpelIgcvg2/p2d9GDHU1NvzXOGdLG7u7q7OA5DjPQgydaJ2BbEYjPlFh5JeLsmSgjKy0u9vD
i7wns5AxjW0UahQq6siPZ3NDD7HYuMogCvjSzKGLMYA9c1/GogiunNxeeu6T/oCgEojgJM5cGnQX
MHE5+LMREPIqMXdBp6ZRYUtYgiIRVKLWIhNG37hdTfSmoRouckanrHiBObwFFAJrzJ5WrihqNf1E
4H2c2tYRIqfpged7fLhG2scGnTro5A5eCCP49ugfUx3HO4RMupydIZ2nl98LLnYhkSA4+eRZcfgL
ydv22UqeKHSgieD38hzBe3njwmlUMyZu8xPB6ltxu/++n/c7sPWJNaJbO3Xv1pS4AQLwxl9bh2Ml
R06eCHJmkZUQDoltlWCof3/dgMviwROR+PKPBVBrd/qOiMYfIUps5UalSyAnMY6aFsClemG5wFJ8
4a3xGp+BtfeCsIfMjEmGlQn1h1LJ0ODqzKf3GfDGTn7X3YQ9iVX2GLCOdI9xQDC3Qit6ZuELFO81
RYeR1NeOFH1v3fQX28B2WqvzT0xMHRQV4bZefpPHUyLXixM8p/g0EkmfPpYEhUnxBt7c/fVz9nM+
BIbKl36T+bzmuJxWV7Dw22eMpU0OxCdgS7z9GuhEETxiJOt1LRlfGLBZYtY3iK3MWotYlSSmFKR8
4y/rKeckYJbpKkrjj3MEW28nPgT3kqUnLkpUoBr8E1FLIvunsnfuEfT/BryLUFKTiG+lhefIKfR2
u2xjh/+c9eyyX2lp9WBpZmiAxCnDSKPvx5BoTewKcnkbJB4N3Nc7kJvsz/YfCIC6eBnGBnEqyPj7
rmHUFiWX9EXIqJ2o1PB3tTU83cIxCSz6rzJabe4ACCtwmisGKTFfbzV4CdHF9xLR6rS8h6BHsI73
ftWSnTTFLqBTarQhlkpJARDoFKhytrcB6YfLaKWPZ7xmVR0qlT+9K7sg7yVpka646lRG4eEbtB6G
iS4+EOLmYaT0OGlSm4hWDdEQAgAqN37FlU3VTebU1CJcP9U8kEYziUQlDpA/WJEeqRyg2OwsIiAU
RngbOdiU/iLMbboRqcH2kyMfvQr0UrLuD6qF4dp4HbHtGYj4nyUcDFrfMmRFw9klMQaGysg125cn
jkyNialydz2Q9NvRE2PXkNi+lLrOXquuEOAvjpdHv8uooz803ewct96SrKSNP+zrZ9PxgTfLz5JD
s3okN+gxjRDadHvbsXxvE7OIQpIUMLW+qdvCvbWsV2bH2xiI3nAgoC6Kk8uLbqtxsotmXIdQ9AZG
bjhdLiNgAC2cZVEjc3s9fwa5rlw0MGcFaQDB0QR3tzoAFSamvyQwKkPnI3R4B0hmmksXLgZrTDu8
2f163TVUBqEJmCxiqSt7iP1fd232V39/MKaXO/ViAOnjWARpAAVxqArL1YLmf8spVEXtxddY3dkV
jnrg3e8iAbRwa1IiNZAW5LwArVilUOYiopxXvsR0/e0GFU1qPnylqrj0HiMB7qdEHRhGok5hlXor
MI72bw+2bI52e0ez39iqVIkbL32UZ39qOF8jd4u5m2jS4NZWmijX1QCBZfnkOf5lSZj4WGkdftlX
bDdkVXLPQfvJvyY6jmywrlRF8gE0X7PNqzOzbjXtRkvyuFE58Jq6YcV0JH7sfYQo7PbWRRy8o6LS
ojGgMv1iAspytoj8ugeUjG8HlN3fsweH8jgUs/T4PA+X3mOeEhF+t3c5tFzcIeFNyipJ8ecXJelQ
trYitmLWZo/lIBhKsFWc00vlOmskalRo8p71jX7fIfP5YmTgwJXpvddci47sBOkE+t+pCuUnWzzS
pySSWfmTkPgDYVq+73oyThvcz28OvoxzhhgSGi4INJhdn/nRbCm01xMtoN/Y33eLStL+UDgCJ8CY
FQGiH0ugG2e6dwfQ2DzUsTsES0LHbxpPfEGXRQMX+XADFnSsm8bnhkKf5JFxNpk9qMDjnjZmEfST
mWN2AA/sLm3c1425hQyGBk4edXS9W5gYBnTBMFkV22t6VqIk04zJLDKcg1lbQPFhqBp8rsucL9O6
xdOtYTZR41F0ZnE2oV6VFm6b3sactnbkeI/furqUpkH+thuftCx1SuK1B9Qo0Cb6mFQxeSPT2IQw
KZ9SYT4Oy4X+982R+fhris98A78fxcQRPXl5hSamtTe+SF1AtL4t3H0+SzfMXRecKz8E0V6rZGcU
QzBt+vGJBOCNZ97xxmLVcBYh3ain7jvuPAjZ4d9+XheHsEQdHaoyZ8ZuwAn4wv+qsztICysJmztW
r3GS9zQJvwz9LKbsySAwOFjAqhVe+CTto9Gvc3xoRbNSCEFdvAsQeIUnVawI4NK51jiSKclKmQYf
IbiawBmXUcDHXe2pQJ9ygPwV/ft0UnspCfBiL9rm98l8GRkh4K4+n/W0sC3xp/S0q2h3rYBRATmC
MmnIc/KC9woK5L2WJKwwVdLKXNcffKup/zR67eTXw8BtGVgBeZLSuJD+PZGWd7VEHXcl120QYW4b
wyapn7zU9I+UFxQfBFBz7HrmmTCjpW3f7vtbpzkBat7Xu4uFJd1z3vu7zjkdOrsPyCwLP5fcu6+5
YP3QOjPDczo9a6pi3Sh9LWyPQNo1WzFOCmu/0UmIx4fjPL5/VeoS4GgGAVfv+PtFUD4OHMUtHjte
BmKoVcHUm9ULEdtGCLoG87q0acHMDeY6LMH/XHaYghaFWRRppu4s4kSeP5aNErylopRoZSDz9sj5
XxweLFJsJHEbKJ/zXtH76zPYLa93lTZgL5XA5pLOXP/undkNBpW64xLnCuqPvY1P/+hJyGT2ykQE
d/Z6yvc0XEDu1MBA3zCrOcoK/lgQCMH51cx818AlAKXrziRFjNHcYUjByH0aw0oSkwbNRWLgcB7y
qlf82y03ec7R6gHQbUIWu8YTmiCm9KyHsj8fEz7xb/pSS9XTVIvgYtqwbtpQRfFTSlI49eKoDMNj
JWQU2d7AXQynVPfu4/Bt8wlJA+maOypX5lfUPIndyDJP+wybcAWpWo3Uk/UqDbyLe+W6cluatIf4
c1zmZoIoA6U39wn9aJJR8YZNN4Usgri7QF4xShsh+sWpExJEW37B+BxS02WKIqVubmCHY1CBCMGF
4JsUI0RG+TLEztGFk2bfElDLAzkvvziTxGYmyDarJL8ZVFcIkHyR67LcL6ZKiyg78ov09TrjmPLG
zz1CsI88FPkVHZqJk7i6NcmcoSpw6OQ9X9RWZNdAvbjTG3WdMhyVsBooiyTecF4zsmuCM2bsCJDR
L35KpZp3uYzPgU+/UvwxjIkmbWrzyAU49nBImR3xP3Zl0uRmCaAVb53r77Wsl7g7zkZJZgAPLrOI
AyHstJ6dFJq872EMCHkVrYt0zmEoZ7OEOAoyEL2Xf4GelBq+KZS/7xLZooaaYdYAM0BpaL1GVfr0
PzmUKRLn/X4TGOjTM+zRXmZjunohg1N2MX9ERgBhusqASEmvapJYGWKD3fWm/1Q4oaIVifFa+V6Z
WnMoQLsTbl5u8CARjjBPtt8MX0MNatg+HaTcMIr2UG6J+ZTNYb2xFCeFP7y2eLmOF3BzLD3EjIbP
i7SnSyatez9k7UjujVUq+EGbovWDY67BCEAtIzB3Gpl7J8L/dZedTYMAggN1Qzw8SaALAzTlqdFo
le4SZGhceZcMJ/u62zxgBEWN+5wCa3dQ72+lv+s/qlgXfYHvdSri2jcoY173O6LxPe+4MkN2bl8K
4cKhH/OTjW4XV8uFSYrc+FvVIi2LHQkOycYrJQ6OCiVMgmb6tlECoWdrY5t7Jnd8pY4R2+PmNbV3
2u9y58rSAq5AJYdRXWO6fmJJ2FZg/bKEdtU3xqiNrx5BoB8PjuGkQHgpRr5VldthWPQtNLVkc4/l
OuwVJLQDRsHlQforVIn3DhdElFFc9pYPgN1n0vCiqPnI7DnK3xihe9Y6JgIVTFkfKnaZCinrUBWK
RwKywRKfmj83buAxuvKYm8btyEokfgZnnd3n11ergnvpIYoWDV8yQy7mlX7m4jzEkpp1PmZMBvE1
nwOd1vD5mOQyxm+W9UjKiroaddCd+rva+J2yw5N8QK2eflg2p+LULWhDCdjfjtkF3uja49+5x3t0
FBx9j5khWAN//2uG6dRixV6XuRC8rwaRi2xY3XEMDcMQviPVnsclxDO3I0tSZfN+80vzaM3GlSJd
0mQpEWzvr43+uLpDKhPvDhuRZjtl1f/rOXV7nCzoIHd1EdDJF/MwHoTIZBsCXkfA66w/9yzq8PF0
FhOHtseNSO1gvnLbH7Jr9mJ3k4ADlEXLbZDiMGVivo4FNcfG0sMl9pPIyes2ZXG6wbENMzqlg9d0
iSLM7WgOzfwlmZNdNbI3u/oczJUTZfwa2Q9fpFdeFpG18BSdmOLDinJDt8RTu8sbF5tIDIquX9wq
BH6UE0Y997LEv1h3MDajbo3jT3YCLkkWs+nN1HWlF+ezbLeH/BRVmCpmMw26Qa0emdTThzNxznw3
YLXjHRQzr9mqpb2xNhNf6hg6PKGYuHjPiV1FYzSpcCKZCasrEnxbmOJmvIdmGBXfjqb4PqAtShJa
gUGJhTR+85kGFWPvZGKCxzPsiT653sE4i3eb49TeAnfITIyora7qPPYVigNFcg8mmxirUqm6cnKP
FPZuvVRREqkaQ3QniKLO1aIbRGtHFNGf0BkN8fIVf0zzGNVARjT00cvMzfAnlsv18Nrg1gfwjqzi
QbqhHu9M/TE/FmV6eQWiQRK9h/FR4qOqgInSdQB8sfI05m/eCJZPrhzJKJ21Cc3SUmiSpBWZBK/R
Qx9lMugB54F11ppKaLLanOZiMpeBpM8K2y9SWpDD+21VcP5iWPEHtDg6OT+6yaFnL5ZD0ZQOaN96
Kl4F79gPAZFQbqVjcCzv5cV3+XAEIIIF9fhIAKQr2NbQkIzHMwiW3IdihJfWh5D24PwfplhGMZhy
fFJN2GxzDX0ud7WWhS6tGmrxx9TVesOLx7mX1ehLIVFRqVaNw9eSRUbortP8CJi1PLBwNUzd8taf
md4vkwMnUnjooRG58BVgrhTyDKbEpxjP9786t2y+PgD2pd2txlWez5oysfrDT8L+jty0JwVjAi1N
JAsGHMAL15NzSLYRw05ZWRngCZWtW+kj6qy2neG67c9gEKDv7H/RJigtl8mf5AXdOf5if0W/IXX9
xWW/13Np+YW9xNVeGq7iHd6MfLJPHivYpeWPoRYC1AMHFuYOPV2oIxu+K/D/J8V0nVAXZBmaDkLr
vBdBmBGYCj/j6DI8+Jxwuj9fm06V0SbUJPeME3Sz26vOUY/hKVkWn/lIT5vx6BXP5yZU7HBVlwjn
jptZgoOvXmxEZzlkbe2Oehbg+XL+i8sWe3Ue8yNgb2nutWJtTYUWE9QnESqUktyPRpwLfoGCfbRa
90/2r7EKBhna69qqoyCt/sP/9qeXYaX9AwYhzR2D63a6pYQ7w4ZZIXWOcjarISATlOog5EXW27cQ
Xez2zA8H5PIfVUbnCi9C2zhwjH15yFT4x/buvttb4+eEllFBi8S8MFCqjepl5UuP/HBJjCOamavy
+e1RSZsFotVRDrA16wDxbQRd4kODfZb4j9RBZ/zswhIGqi8VAjg9lYjlPQBr8O0maJnxXbzv2T2b
IYlcnoLUEbDjl1N4pTG2tNwSxSUVmvov84HbGYgI/nahvtMxagPCPGiWkWyEpAm5/0ni2ULJlewv
v3aY8cR8s/Y9Ec6+GLYN5K7FpqrSQZa0qSuMPodmHMpjAmSVOfy0zHY5HqdM7IEcg6wYVXB5KqKn
OizNb083MCl8UY4VdXNV0tdbh9Yo6ek08Jzyhk8r0G78QJHsoivLicgekmNfQC5OBUfOtAqyVqEe
oM8IHKS4mZEEBmrs0+/IZu7GHRAldLbvD+JRjmhyDCVXFgetZ10AK76PAPt1oaG6nv8fURbUG5G4
hDFjvPVMqSSG3vpOA5Tq7gYDVarzJ9lnw/8e5VUgvDSiVWLTNgpmlHEKklXAC+jK/t2HjEwEi+yI
1d8s7YUAlutjvSdxWsnL8EOWPoTf0kk0PAOhgAWwOealPwGW/78v9Um0NUnzadl7ulsUXIrs/lZo
CZ+gMUM+u2Swcq/qcmZEh82xgIc/P+WH8hYkuqlADshdqxKGeJfZYpQxmoE/+yM5iVJtsWXXw32E
1BV3GAKguMhZquYDYcLLKBvAFhw/JD+nsZT4ZedjLe6Z5+uAWqSPrecIO8v2Vjqt3NmOIIrV6dn2
lhBWOGb3pnuX50ME/NX0xNsacMqelZq6DpOWLuLHEt2sO/lRACqwh9m35a2s2vR1QN5ERgniIgNz
jGvdRryXDjQi7GW8CZWlb5mnQVRka0Nnxp67a+ilCD42J/54xs2E6Cs6wTRkBGncGyEZ/0aOvwsx
iwWKLNd2HzgwmJa1cGTZaq0uf8de8BkTnqfcTqKsjzOKRj2Fgjm4jtwfIOC5rAuJDIimEUGo1ssu
LjxWlv9yLZM/Gu1+H+DOo/7JmcUhmw6BKsfEcs8Y3ohtf/ocrO8W8lS/v6HieTudMfXIMs2qZnTY
lvimI/KMs6X41laQFJinj9l2hr6uaTWie56MtkqSeicKfnnrURNiYOixadkWvRjMfJvk61iYIdfy
vJGx7ocLo5BGlcrQUM4tSkW73S1XHetBU8+1VrvsHflvGE0EPmBYCwDM4YJP48IoQpMZHkpKcdDK
hDduV6WCLgmiUWmLk+KpGeYLuRJNm/kfXIOmGH7k/Oq4uVi02A4d7DiDlfRnd1Rmr2I1QUHysx9s
X7y5/BUpjufj/QTllALvb2iLxUO5U+NFcdBdoqfLbUd1QwKjAq1+vmPCAQCogib321TXIWO+03nq
BjzsfBLWUx+ANflRpJGCZD8v28BJE9IuDuPcGkHBvHxvOGx622YWM9OgOHBTTcw/DBuJRbpc3lVZ
W4lUDUYEUIn9UrYy1Pzpov4g287oWAE2eD5C97Dg8vqdLnDIo/1JpoVa8F/mre/aXyZ7ZcJVRd5M
r/0sml8O4YiBAZ/bRQD4p+uxw8+CPB5XbkwTvAjZezOk1IeNmWbyPc0CtjTzZKf2DYlTrxmWtVWB
JzZcmFu06GVvGNmOfBeauPwcyNhXtBJ5+owXKpdOZ9Sk16EWpq8jPWwLT/UKeRK1QuVOlTkO78tS
y8KtpkZ9b4LMvOval1rgg7tK5f68044DpSOv9bxdpXsMwOPzfgPFdEbfZR9HvYN7WTyZhkcFBV4j
Rmv5SQVULIZx9fTbTSIsTAj7ucUID2OPHc9g/jxLzOrTyrFLqiBXkZOk9+JFLVMTi1YBFbzA5Beg
3tNsUioWQvDTbg557d24Dh48plhAb0/yCtd6Rl6sC73Nxro/6/Eogtz4lNhg9Rkyj2kpTbrQJjE6
9Ol+hq9Zt90++RvpOAvyFVdBQsZAXqbjDamBItUNTvNLOkq7rmR16e4/w2pk1/Y9LB0Xz8nMOy/B
QOwle0/tOOUcwKhx+OBWoF/ORn8xaWkWAAZHUZA76p8swgPTkvjXP6RTfFvIPpEJ7jsDiHW9ZHbe
SE5O3OlJXzGWn1wlzFa63NZioLggI+k88oN2hYL9JZxUkLtpebLdxNtJk3PiXv8Y8amwVjkoKecQ
fCNsSZ3kvS+XWWjf1Oscc5kDTnrFi7XajEwglEvfsezrpV4WR5T1keiqFU1iTz66jmlDmpy7ZyLH
mnkyss5hVB8pWMWfH+xEeQdvhwiPbC0h/ufDHfaKE9VQctv8nrGPVsnTKYOoZo1pRbWG5oaBZthT
nqr5Yz1iJTPPv6M8uUZh6u5YTvVKr2LZt2cJTM7anyn0YMbGs9X+T3hV5Kol8MkLIibVItGCU/GU
lWtxOpq36IUI5wq+VD8LjJIjAQCPokqK752mCkGVsn517B8bpiWj66I+cp/Wrz0I22+O4Bz3eAxU
1Huem+yhmlYhPuHZmcPMNw2nZWLnkX5Vhc30ArDbKe5S6zyHU4hMtJJvJheDEDS5frCOB7ttvY7A
vpwJrlHUjsT+fc7/E0uNXVYTS51HTuXoYTX7Qrzh7krruD4A7qdBv/rLDZXioPSCfnZ6Q43yD0pl
aHFYpbeWg+x1eEANmeii1WP5PqAH7GIZRgrsG6waikfezQ0XmUoiQyYLII0eR5ux3o5KUEDkCusU
Xz9zrCuWAu+JPaw32WdZinYyIEZC2bdjqI382vFmxGztUkyL6bv49DXE+qvukMijAlXdrOR+un6G
Ac1ACun9qMvmsk8qKw1A8NnD4GAcZjRYn8Snikc1Ne7IW99zIT8KN5Zw7r7KQc1sPKwN+UtK2jgk
Uk6e6TXSN2yPRDVdtxVAZl1dTuqcYDtUro0LomoxjM1SqQDnLvmt3EzahelJNFQE1JwqPtvijv4v
rEfiK0z6ZsPqJBhzPEdhE3rZ8+I+jRnea7AONrE3QjR1f0kujmOFdRF100r5/P0i0sLocPC5ZFST
+KchPov7D2t/IemB53pBF/9mv++9f0s7bWqy1dkB2/5/gZoiQ8e1UBrBM3TxxRq5dOQhrIN1f5Ho
dgnYIwSFac0C6YqLFPUUHSYZYCITv5HCrzZZjEuSaHZPEkqXxnwXTMBT+rIFl5FdijyvlMRk2eAH
NlYNIcQ7T1i/DI5jl7WvPbwIYbmvMuooxPR++e7loTpDcvIe4leS+s37ppnALG3FAIW64Yv2ZSwp
/i8NTnB4viEGBoNWeKM++7kD9C3PNbnnTiBARqvVD9BHeW2Yt5vvuslxNMpK21wMaQIirPhn2ViX
JZGqEtx7u7BVc7ecuSNBiZ7NiHWkTYDdF6jcYooDAbc4FJfNwwMdPoVOAgjuXo12BueyKrDczWRn
S6wT6uYYJi90vynchzMPo0Fm/3cOBuuJoX19fb0squD+7KN99xDcdh4/7jegzVpeiasTgi2gP282
grLEELbwvUtR/MtxjeHwl46mBmCoCS2NLjsYncGBN3kELLFCmd0ucYRwzSglbqN9sPazZz+L5SDG
yaalzw/mCxoUiLb1AkeTtjGipdZ9k4V7YRDXf4hVnlwfELyQChsIJGaeB8IZES59aWbI98ZY/V/R
gcwrPgfc1faSnZjaxNXPFDBNTd1jiYTpbZCs4qV4p+L4uS6td8pYU5AnTF++v5Co+cSpfdsoOSaU
BQJw5rNvqB8PFRwcNgf+N5A6GmAYDQs/nOyNAvIwlQqHq6zgkL8BR3E8t7qsoXfK3IUadowXI26P
qtlj+rF8/afqS5oTNTZugbicWPTA5zD/OWJRTIcAMupwSRlqtr9UZ949Ia6f77QajQatLu0IWJS1
zjlSRkiCBm9LyLfPZcQlI1fowMqe4Z6ldKOi8UHSE6jiW6kbN+MDe3DHiDwgU32ndOmpXPrsbwIP
2uR1mT4t/EkqTESb+tCczy092MhHzZkMw4jZzIeOj6AoWums/iGN6Jr/G2CLmNhuqOdSHvHTCsxp
Zk5/Jg5k2i1uzbBYxVg/eKPTWjwLR4sW3gvAD+JLIHu9s597WgnPpjS4A6L1EYzTTTRNHaDFvlm6
AjnY3vX6nPVa/Vn7FcYFTmIRWQByfp7TqMHCfoQ944snmMqVXDNaNJvQpRbP65EEPs4D1KOSiSyn
KgUfnfByrcCeQZoo8Bf3TfN8BrkDHEGyfLJTyl6l6oxGFOvamtj/2dlmjakwgoqkZHeZTr4E6WqA
ePQTL5Qg87SHfEvB8zm8faEhLmUqqr6AV++Kki+PUP+ZHZ0AZOo1ll4WiePDwlSsxijyFur31J22
sx6wTIuTUMC8q9xrmScn8Pi8d/6+xvhaXR8Dc/Qno76zQs8KjA89xF06JfNsN5O00uX/Z5vgauNV
RsmYAnSJlZviBdPRohEojzVHpdeakGijzyVzM1KkgXHsspI7dseNbftNzuPc4Z9M1749lY2U2jyg
5uMecEFUEHlYg6XiGdC3AGXCCvWx576v+ESOgmKXGyrwKwLOqE6DiwXwohZtr93TEfNeUXhHAyYo
lWfrXvZH1q7wFbynMiJCgJBfQ6tqtOZL7gZaKFx3afqHrWzXI6IgGhA1kTKbU+AGJfiWUWm4t7Fj
GbQGA1XpO63SYh5nvoBbXsi6cMopk1NojFFLKai2PxzhKqpBiok9HC8be1NRomwRUJDvUWxkfEv9
lQ37/Y8JH7Ojz26f+eXomB/kCbp9LXOu+GOTCD7jjxLDoNaYsclrjSCiLXcuWT+NlC1HaPqrJE08
Gy+WT1E6PxeYWhUDrdBXd8nQBc9jXXcRMUb+3oxRIYTmJn1AkEsE1tfVhsJ8dCvkwDCT814kXKmW
zNFq0a8BFeS5nIIREPcmE93y1LSlvl8ty397JA4MKGNxxXHKONgLL/aqMbA5tfoMi37PG1OYwD88
Kz59CvxbQkuZApks/JmZAl2FAv8ngSWhgina6mnyY8tGXaTptYshXXQIv8wRf5g3wyRdPRPGTdmJ
1qAUHew0LIs8FzJL2rlPp3XZwem78mkM4pT45ZmkHBBZTyS1XZic5MO3FO4JkRdR9ZtJ8/9+a7/1
ot/POeBpO2B0O6uIeU2NA4zmRGIjxe3lGFPsTSws3p6LYllPCMdVrbAh1OMCgaedM1yurnQvo8ko
gN504m6YVEtMyzo8MNdz+ut6MH/lOxpBK9ObyihURWzgW3C7NaiSW2WBABunUD9rlDl/R/ccEI+H
1Dho6A06IPGTRCGdNR/Rq0VbiyBruT4RY8qYj5qL+AdyyCLAVCVAa97RhL0FjQAhFKtSzo5BEYyi
JsJRYblQKz6AV8VMKvO1YQWnHmKUWoIj+M3+fefs0/lPqRUVvYVHzv17oErr8k771n6co2jjE/Nb
owo0Ge9TYCMt3P/mTN6RKQZpvGp8jf9oWPGgvAAFBPhkFqjrgKykafmnEZc1EIssoXKu5DnAFfgH
lNfgJ3NTxKVi0SzJuQV1xvD8pO9hx5IHEN9ZoG6UZBu8aWZmTet6k9QkZQr4v8RIQgVUNhwKtF9/
n4YIzKiLdllXeqQ7O8IL2G3aYMeJW/ykKejFund3mGU2HaAYkoBwOtmIatihXb+jzKyZr+0o1dhI
nZDn+dqqznbvyvEBDIshc47DhLrACKoXFcgU6LG2fNR5CFvJ4IqCOygIO1dZwxDZltZvrvw5juCw
MQ7oF+IBxoBq/gPsEHdZdik1SRIRXKSb3QViF8TGSR9oqg14Yep3nEosUsDlhG0pA4K38jKKck/h
qgcJXlt7Ku53lS4LDUnnDKaVMbTgFY3qGmURHCyip+3rV3SEoViJPnptQQnkBLm4zeIGeEVs+FBz
/dAWocRUmkkB2LDJfufcCDYw/o05bLJvpoDQ38RtrwslEOuMstW/Rx8sqUHJ+0g2glGa9nQxmbkn
svrGB/vPdmjfm4+AyGcw4ZdLeEHmbsUDmsHWISCHjPf8FAuXkpP6YwfMLrexjORvxpRSdbvh4n6s
PQRElA9gBN6Sb5XxcBM/TyIqaz/ixOHwwfXs4jDSKq5F8PK4rtLj9Vvw2WHUJjIF3FXH3tUKXmlZ
ZuBenMGz+TjfqM6dKCUKCISFau6zCcnNnBv1iJDMWLwTEWGpxz9P8KqDe9djg4Qg+NNQPryx3Ot9
AtL4a706W4EaV3EZV6kErFocEUqCzdFIICONGZOZ4Jutewzok4L9vCy/f6jfoYEbBjHJ4BpQ2s2l
v3oKYqOG7u0tFOXSWmRS2fLI+EKYfYpAl5K9AKggs2jquiUFU3SzGD0je1NKdWxIdowBhJd+4Jit
NgcGFORBT2BF/O+jpXQ+4RiiPnAwcoTsCHKgq5cckHdvEAgVarhuV6FSdHB1xOgcClxMiMmZ9l31
1KHVW/D/MaHCHp2IFj3f1Pqxl+ABDwOltBuNt1kaEmmuhHwLK1YWwR82TBVNtAs7mNYNH6ZoERbA
v8k+OHwlqGxFlJufg0hPFij8jRlm0fTyyIja6Jfan24ikUFRuTRHZJs2EbHyOEW2qgaGv/uQX1IN
FJTfqHXPGGFEC04t49O8QtT/9mngAXVt8bS3gNqzKboGVwE9dXYRlP/qmVEcDFQRzTPkPst/X4M/
2y58ESwgB/4/yDdfTjgnWAmx6Lb+xd8yVg2+ku3BvJ5iFjCTtCx/iF85DSmqyMywYpRvOzHEd0Uu
GYuv62S5M+8C3wIIi0KC+ZQB8oSc61U0ZhcFCAHbVCWz0csYGVgeTmhKcvUuRlt0I+hThXnJSN1U
qme2FXgtLtENgLJL9EwXhgk3BtYB/QWUECJT6BqVc+bwAr9EQwl8lBBZllaMHcfrxhlBg2lAFkSq
8yCX1CVs3PNvO2hfdirDEdRiVEQdU81sZBl/03Z3o6KBBpUyLkY3xd0joy9MW3I8NrAyLG05AUqE
HnAN0WlgBCDs3wzWjsS7rJCH7axXz2jvgirBRP5dUKMimiYAywS7DVTQjK7eddX36xQJ/ElMunPJ
XyzUnqWEXGt/UG0kpNGP9b/T75YwHk2ti65bhnWYraHqqx/5DELw82+/UcXXNzFmWAFf++8iCY1O
CXLMV7n/U0eqz4m9UYad9k2ZLwg47akk88mbb6M2/qDtRalofBeXJ9SN+OQN5ODsSuJ2P48BJHOK
yqENLvKeus6BPwr6Sz1+6f5mGtEjtNAbj6morSx9mPpyab6iY22+OPqyqO2RNO8caf861vbvxfji
Odw0LdOowL+HyFC39rs22vtNU2KRMPrRwfbztiz4zl46ir/n+t1yV++k6yFj7+zryBgA4MQRpsml
yCv0XO6jeZGOTaTmizuQ/fOF+z1eRYoioZ3csCTsggBOQn2BFou+MBSNQ9V3WZimkQR0hPe5C9S3
w9D7X/lx30kcT52U7qjQC6kYenKSCDzeWcgjlMaLoPtF+FGf1Z0zgRpYyl+BGcTVZ4TcYxO1XeTU
EREzXAnlj4BP/9Py1oRDbk2/wucMv4wY7tMLhS7lC3kA9dmZf4kw1irUg857iXa6+d5a/mdaTMQT
zBxchk2nw01ZnPI7UW9vHb/oxpIGOo6HgHetzNAgmixFGFljdzkavyMQlj0yR6AHbjNNx+aW8Ld/
kMVioY9kF0/l2kCUU00/KRwpViu8IpMW6Um4IQX0Xguezz8ndH4owZfWBGU9x0sRrIaBr4BxN/C8
9SXsyWVeibR6Fl4DG5nPZcGvbldNrKJyBciP24wAnq5lVsn7xsiHPZ8y1/lNIN52PGm58BrBCjTn
a5E3jIX5T90Tu3PxAF8IRK+rzRRR6yBV0ZAIR1U472Xy+3QkDyhXiECFyHjhl/bqkBR0tBWYmFTf
O6/7K0upMo3vmKesZ/7Teiq8WOeZ3c9XfEooZYSut8aaApaLZBdYFmVbTGsevbyvTDwzGKyWOycU
xIl/fgQge0cBtWQCc0VZ2dUTEsJqHY9xH7tVQcb+NHz2A34RuM01XWteeD/LqVcRsC86P/InCybf
MIgdfBDrCdjZBe3+Hj6mLO5dKch8ktJmBKvgF6+9VNRk0pDDbfulE1jKmlfQNOGu5/OGgxDfU3Cp
jCOGDt58B10K+fyTQWxR2X8MuiC67d8CHylBVfiAv2SXTx0cV34YxFt2f3MpdtwDIVFBvsmt9Jn9
66JSgGkSUPwZDDCLZtuBLs9Sp1UuAZLGNzZnXEku86SFFI6vgRWaBoyRCg4RlR3V56pK2kOQ9OV5
rTKiqKTC0SDOPZbv2/1rYy2+EgjIuMEuDy+Q+SAg09FFkUVUC5YvUX19AQn1d0MdGsURR6DHu4nU
yf4QBj9ZaummtixiU0lsqStlFBef1z/Xqpn8qWGSjT7uvPLPd8oYtxwifHZtpWkDVm/IWIthvQUM
j44zroiMqX2xjgM916bUEBCKAOOZFMx3dLvEyjP/qZqmkRkCuL9J3qJ4Ky+PMoHS5uvYJS2u3SW9
358cWDXM8CojiMC2nEcPz3bxxb4xUQx1iU4AdFBlzsR+SOIHTdSR1GnZMYM9XWWTnVLOM7xbD7GI
yai/9PoePWEcGN8w852rjqtPfacrPePnhOiCz8bLzGY/sxLD7itHCUoiFjFGyKy0JIezQGJnbof5
2AbaEyq1sqAAgJ2vvJsHER81WV81KHIgy9gaXueIz3rn+z4sMRcWRomuQujgoekZo3+dWUqhTndh
dK2wtqS26YzUr1AO2mGkiCwgio5Fd8lr3/0oue8tEBHaeQiAE8ITMawuzS2NO8YqPiBV1MH1Lxp3
RSFMV8cHsAgJcMLJvn32jEImJsfySv9MKFa41jOSYVE3Bg8hQoAPZ9XRiI7gNLgcusj9InPoTuhq
DkQ3lDGwIAP/iv0O3+1A03BxBrGuXLDGX1xrsOT0wvQBVtMezFVTtGjS2gHzpJDuYC3XxeXMpr9f
9YhrRMX9lhfmzI7sE36iVjY3EsWCYl5Dz/kw0Htsl8uO4XsmaK1M5fuU0Ga9dslDAJhEoIizer9z
LqotkNX8psWD889CIzxECzdFUCHN6cUKJR+J7CDkAO7wRARnZBPyegnQIrsmii0lGKT1RM4pRM+h
MPUVJ+UlsC6ujxeSHCsMjtmcTy3icU/i/Al+RQeCSaOw2cjYYWMmvyYaa/EnbD5atnUVR5pkQBBx
G6VnbzQBjwYGGZBqBttr/BRqaPixkNLcQna+GdAXWeg6Tq65+u9/sVN3CeMnXqajZHOdlSB1SJCj
6uBnxmDtFyNEL0d3U0yTtVUFGh9PZyr9WASqBuI8bk76aFuBRJBnKxilGVysU4tQfI2OlqjFfbZc
w2TnYa65c9O11NKF+Zw+PfW0HaFR2IGJ2Goy43GLHMMUx0q42lnW02neY2To3/KWAzeHqaDtd905
m2qSN5bYQ/UBeaIwkdHRmF84SEANpkuxgwYj48aVAcEQbP5+vEJ3w+WiYGSBU2FEMPRpmR9B6ec3
WYojCfWPAXRDBqbdfRgsXOrkQ4Ebsb/ocZBRmbvJ24gioSae6GX5nkKYKNi0pP7bngH8REHiQpG/
2lRuF3BT6Ktp9S0buuQW3Dk7qSSigPPv5wKJylYUf0y/wbRblc6XHiXthAfjW8vsgNT+vnnv25Ro
/1TV9sVLJrgcicU4tC238Kb5gE+dJwgdAAzKVc1V8Hb647T5xRwET2qubbVVJhJf20+ZKv1QOJbB
zdPIllg5NuPJxS/OwJkpd4NY7l5SuUdnhQ3LCfHYsJeuhWq56wqIr97EbSl3PSxfkwq1wgaeXv++
TujXRYWQvg4AlSyImRyj6pLnBPs6ig++UsmmOIZEAv/yDkwVxQ4ldlbFI/3+40MRbLK3w83wAAQi
bN5p/r32C9NuQN9gri8S0pE6ZlCiFLYV1JVHsucjaxS+fSykueY+sHhC4XNBlEgzsByuC6w2X+Ik
GDMFZCBf58eCe7rWvSdZXoW/5FlhGdP1vemwMbACsln11mpZaTI0kfP/aSIfL6hShEMqmS8Ph2Oa
uXQeOUPylhxSCyOXadOLo1BdCpvQVaCsprw2pNmFuGjqvBYZelovoepHkiRkUyjxrQWPCtEkOrTU
QIBS4VBI3MXXeFAVGlnAMUpkz87dUaYLWmSNme8b/Rhdy5Q088DJE8m5mpwtS+EqCygdeb6hlM9v
d0xQRaDnlDjZZT3FmVrS2xow64UknTSFZ8x9ECSdbEpCzgB5zzDuK7mqg20nbqVxCeLMj1B4DxXF
I9AoUQKXRlrfnNKjThcr5XrUK65fBHiWN+HnVoeQmenJzCWBM+n1jfIF+5tc6H6d2Xc5Hh0OPzIA
A23LFRnBX2/xD1z6pmEKqJUkiS/nLsZEyUTcM+sv/rn5aodFu2RDY3xXq0vjikcbqMDkM3flsQ5u
6HpfqEC5+Ip9+VBiYTtts6Dz8DiJNBK9ziRcSt3IVNIHxi7wwnipSSS39uiYzJZIVXy9rPiK/y+F
ddFzt3Ke/DHn7RPvEu0z9tynFv+LrIGkAjz5edZBvChq+HG3ttvkwtVLeZz15bQURvHmivShCSc6
n27RJSyfYEdqCEIN/qXvoSbBxyRchwVx8XGj5Qb5NOq4AcTnByuGERZmtY4EusHaLd/atvOYmh+J
nrwqNslszwULwyZNgVPCilFvUIBDSceFV8NPRIMWugpWSoyvNGGSeVEZuB6Qp7EGxP3rHLwAtzOb
m/JTS/0SB8ouc5Y40tEQcg2+4vt8TZX5KvG1dBDTAbQa1HxDiXc7odP0FPV/ATI/lWc4Ik2Gdmbm
C7EORFwNIpxROb1Wcwrda6rxUNtRDt9QC4ja4oDQxVIMpLiGwKIpnHbnpAxnLUJjG4Q9Ff9VqDy3
gigPuVqSqz7ugnQZYwgmQXAeYdsg3ScsqM3GBa3JPj3Ie/9940+xsergOWthDf9p1dhei52PXFVF
Rm2swiA+hPmT4P+EeA+0NgiSCypXtkic4j7U6FBpS/AoulTmA3pMYIFanAJWDyh/uNUnPlR2eIbr
Cr0RYawN+bEfVmWaZNxmDFOrVY7GLPWalp4/2ig3+zI7BEQum9dHVkL3NvEgKkr5qKjPt20GqAdm
NHlFBcZeKJGygg/sy/aJsCzzfOyk7sz3RAhUp0ugYSrNjqC/TBmZ7fzbk+j+ZXoJbQbG0SynenJO
gBA8aBqbjNqjkqvOizfuMHAUQTr+ri1guIskFh8jnKU/T3S0ctKPbksrXdzh+hV9Vb0jrCBVuVCB
MjGh/mgFL0ZBQWYcIBDPS+bt6ZlVrjGzGR/4N73XziDuIxMsZk7Zd9090PojZC5j59NqdRElvJFy
9RK//h5bqja75QVhdW/Nj+DNYG//OtvaUre5COOnqyFbJoFBQx1Chjq2JWhu9ZuDDzRjWMjny3GZ
RQs139a4xQHCuLJqD9hiHqWcV5Ja4iCIh6NwXin0ti5Gz5a9Cs4s6eOP7q16komsu7pCh8IOriG5
Ihl/mfLeGkDotr+XZu4cMOT5g0UKRlRKBNsPfx0JmbqDXP/obF+N7QkIfkvFvwaxXX57cZRyPCbl
l9AgCbrJ1LJdtykIPz9qorL0Yxxa++Us86iQaKBKQ6U6COHeFJnE/xBYaBaMeigRt35/WT+AbQKo
jSgYRWXSQqJOt4RaE2OwxSVHNkmNclSjPaMsuiJmFZGp2ic0bvqilLMO+3Ts69nDJU0MLrfzVt6j
ZHvfp3pSFrmaUSBoaxb1+3Je/EJKiYVkWf2qY7SYDLmMKWhwis4Ina95orBsXvrHpQiqf9kVIjlz
TB4x8RCQ/rpTnxMPp8J2CpnuNJM1W6392GrPOtVNqnBhQ4t5bvXhe8TrmnlR9JvdGfxNT7qsIRd2
BraLmW7Cv7a7s2ZKDcQxYynHjd+Rxy2L0csCQdaJiDxTJh5RkBuXPXPuy39ZEAG8jcGm9Kpb5hUg
nNbzcgWj0eYNA9OtcCEqHKn/vE0UX8SaGUQcfub7Dtbbr0DQukpuBTIZBovLEui34Cx1aXv9ONUr
U4zjqhjDJ5U9ozfsyjmB8ceAkRXMkXweqYm/bwW6Eh8Apk6affETYeoea65XLAEhTprJbcEFHspx
WGWmiEoxnIjfmAxUCVUV4qCwlsujHMmzZj+CCKus+YwokTL6bs0yRE+lu6iBxSGUV2fY4LQNfa+E
owPLdUODPerVwOXzIy/JXNsQvGN8B18dH5nX86ndUWRkrYfDnabFG/Pg52adp9iBaeJnGUnOJKvh
/2FkL58LdAKs+HF22hB5Q19QNrQH6vSDOlXMrgrWoxCzlVaIaq95rWQ1/VQ3webTQrgd+8oltQtX
RP2uR92G7vRvhuC4EzDaC8InkPo8lRMYuVSyrGKVZS7SM5YsEYx07rwRFndUnLJebYoE0Nu6IG2K
wyRWz1Gk34iJezrvJsnrGFux/5i/A2Imvsgycze3+C3Bzc0E3NHUqJg9K2UHyN9kpD76SYYQ4Nd4
+Xqq/k4L//6BrIN5iZFwHmkJn/N5uA6nR/WqPmeWeHaNP4wGPNEu7ltaKoWYlSuWJUVdDNGuy2XZ
SfOzwtKY6yZuZ3T7kjsO0oee/y2l8NPhxXYncLiOQGKG+r+SIg12kpsMuINfXVMv7pKIZ4wk6GTw
ieMqTs+AAcfjhRi+qwmjz/KE5lSN2DWCdQZ5jS7HFfg34WiAdiusnrE22MW1LUu5yw9cZb1ZDOmC
+KGn0aHecmPggE85xviNYhLWyg2r+lwMQNh1v3iDh/bOAnTBgU/m6f73WArr/A+IzBNgXtKn3hll
2+BWofSMBgSrFK3ixtR07nrJEH50sIUPsPL5gtnzzO21suOy/+BMKGP4MibTU5pVs74ADa5Sw7UU
W6bCG4jcbZuvP1WI7YPuR7PuapfnB31wMYTRqMym/U/+Qd9ccskGItIgwrC20pHP5q6fktszJYRm
P5eg51VOvPm6iYw1gYFL5xYDeh8LV/l1wVf8MSDi97DrkHYcFW00YXjRy4OLPg9SC7/5Lsmn7uVE
J6oe0J4jrFQPQ+QRsh7UL0CAFb1V7BxZE4wBxFpZXbXxSCR39juYs136mTORq/CkTLEM9SyXZucA
YlektN9YQiDrawOnWf99j4memI8qBU45JOlKKvPZOGhJ2itrwNOExECn6Hj76ozH8v9ay3R+pjGP
uyYkM7yGo3xHQ+1/ifbkzza4Vfs3mMemITr7dcVkdoSx15bYP9c/vV0Vo60H8gEFnDEaQhpMeJtO
MO6caq7gJYA1kHtb7tBDW2BGakvljAhBvwComovYOLLnwtQgwYb1gYNM9TT4FV9PRWOonaP5RQT6
v09I4HFUDgeabR3SA+3yS7Qy7Ht5coLaiDQuy2NNAQYg1RGtuhOjg444m1s1N3ifj9SmX4Dl5okT
N2SI0dM/gR9eDryQUgcrOnDVChjDBmMgXOTNDoq7Hwi7csoZgFV2yeinl7JIAeXMZ1uG834UWXjP
GkyPVP4edZKpr2VFeIOTL90udDm1Iv+bPpF6HEi7VjBv1ic8HkX2tBJaTtMRCStB7zSVXGDrhe0s
eiXsdtDM9XL8OEeBILm3RRAJWH91L55CfOH3lJQo0Ajsz+d4iqTEIygE5rNlk13JvwyuUNOXfBIv
OslgKKWIUpTGhA2K0QWw5BTYXidKZcmWxVKExi2UK/RxU4rz8rNxJ/6zRgPmaSK+ULvDHB3E5tkI
eStEbofJ9BGkPzLxprYUYBno01US5KZPTmfalAQR2UueXs1J6qh8uyKitvv1upa7KJ6PtEfzL1Vd
c0mywgQrgM6gUbDU2sBi/WpCcOO0u5E7ZOt+D09N3tqZVv1OfEZLPbvpuVYXtFSUn/dQIOuOcOKu
wT8aXxenKcfdmc/1tfpiG8hQT5M64p1PmMLg7WZdgUEir+pRZeSuGL/SgTzctR2u21kjKvmypqxS
q/0aBxmIm9tPPTXH7h7TCGMkNo+0kIbWR3gjk8kU31GYH/pzUY8e69JC93tSMN0HwtnlC/tFMOJ7
2+mS8pSGQZ1W7+D2koR6ii3Pr4Sm6CX08qwn/JObFzk2ezEL81tdzPrcH8Npy4x80rORTFLSlceM
uUSnwA+OPNPPFVKhtWlk++1ZUGO5l55UN4hilkzU1b7hy0zazIuMVfRv5oXKwng9Mz6RYt+2nz3L
4dokQb1nDAaSeFDOVYecCoD9I/OroEpW0jYRPb37uQ63kKkJUwa3fxtnzLVfOJTiCRA2pWqPgQcC
5UWl5Wzd1Pt4rMTUUZDP5FezeBxKO3gN7YEnVxJH7MHTfGEDhUD0HSdCFfxMdAFhJeZ8M9/+xGBA
MhQkSpj87nmx/Kpt9nkRqNAJ4G935JXG68DJJouHk77uQzwFjtA5BPCL4ojwyZ08D5e/qkskwf6w
I+0ae1HAHAYoq3n7ReKeZbsJXq3utrsK+d/68ZXToCCrGz1UxhEIbnFWNsOu30fwxGtUrQ1Cx0Rc
yJrrBZl/Nq5skH8mZwDVRKG7egMRRheQ+Pli35dP30EWBzzDqqtrPOAX1+lZN3jx+6/7OmRb9LrH
a8KPByJRBG++JtHMsQUzBuhAFVnxqbaXoscqonpVTJACiroOzxeY8wSw25cId1RxigICAMW6/yAw
qDOuC9DvLaVHnqoGqW2q3AjapLrF+PXmCGHeGNBAkuL9u5wl+WT57ys+OTIdSKiY78eBOQUgvKgK
vTqTg4L6cQfC+Eh8EIJ3wwXQ9kifXGREFAi97indFFMc8m5qGlhOqELom/8kYbibXLALiIP0tM6w
/GuEPbLb0OjAbvcA59OBBl9piqRAmTs+Jm7JqtoeK+urQR9n7b/JmurJIseI7fJWHp+E1EjxpBJI
AeRxw2x2mxaTncGifmkAOlgzqYtqNsuPpT96qPgBKtwuu7c0bNRIBgl58RJrl4gmJa1e7bsbPmuU
LgmPKc385uGvahfwcPoPC3WJdHoI32zu3ydwos7+7/sc2WI4JzgB7v/0cNUweN8dlPbfBE+OBTk0
e5enKH7Kex5L98+CiR0T6JaM2wBJtdwvrdO+m7N4s7/dSJF1cx/D47fcv+Cx9JP6MfTSSnUsKhBT
1FxU8Oa8sL5Hmjccnphlxz4eGyRvAmMc+Dzi9VFsR+DcmVggrk0BfKz3kck4lHD6QTb3yAYH3bTN
jRrHQOjuRrbzZtJ9qApvseno5Z3fnFU0qtLmSkzfD35ZdaPs25SMc61r/XDJw1MkhxUCGLivyThx
nuNs0f25NXBEQ6TSRTVI88BZqSzck4lEVswgIY5NjJmRf34YY1NoklIFjtKIPpRTCtApyw4ZrmO5
vbRco90Nc2vk/gTxdt5EUJon2mILosA6RLEGjjsUZYvOAR14NDrwjqE81Dh8nBCj6ou8BPsmWKqX
z+RwNqZkNz8tgEVIqCPLOaRdCI6ZeC6Kljd8yrbyRL7hLTJTuDsxz6uwwBuoz1GVF6/Hg6zfmxOs
mV+E4My9ioy1rYC/DatiB4MwLoS8lgfR854pLar6udILqCgUsqNWrho7gYgSTpsxEeMMX4Hlb3dy
V2Mg2g+xtpCR8WWe2Q87Baraw+EKM1xOr2JRluxCgVVNN0TJQh5KN2+vGGQLWm0/xc4GiQ41ZPLf
a4tJ/X6etAPCK7IQRwpsMJkeV69ILUE9dPMa0p1LID+yyPagD50YgzRP+pzN++YY6zU2aQfvxld6
MGaPjbEHSzTEBl9qeptFbTInN02s4st5FdcwXicbhsSZ+b4+arxmZbNPdYsrIEpK0Ty4zIKL2txm
xvnkTXCsbkzhcALhHdmKrbK/venyA9jLwNhOnPgOhBwiaKigtOpEEN/gWG7O8dvxrcJ/GlymWhQL
i6FT3kby1DjtPtCGUGaL8ru3scWfMVSLOrYPj2ozmfZ+SknjMwRI902FJD+KatosYEdlZiYWSXGy
hP33iG9cv6AOJU41LSnoLxb/BrOvwy5UOsHtEyYZo0d9j9vbR7X4yKYC0lqHcR8ZdKyUhqxMR7xI
D6yH/b1Tx+qyYxW1xzl0czebCO8LS2YD7C0xqyKtLuiFpaPZ6IVceaqlchkzb6KNLw/DKop+c0nM
76EQnby4mzw+Xuw9avpvdIQpar0ywlXgQn9PvH4reQVqaA/n5yrIGMuHVwGaV1Y/rPXuKI0O5q8A
THxaNAdYypXv6hXAT1B/7nA4CDw6O2ORKaRM7gc1WSQVDnXR22KRSptYIbFVuZuiNESKw1IXkP1G
Fxz/4+iNi3d9eHxKhTJkkZN7kl8eXHKK4/bKxnwbRIv/8RHfr7C/2JXCO1aPG2moUE68kVArnL98
TtQg80lxWK+CqyQozLqGQPVrBEoebmWj5Oy47YOQnafQM0MW+9E+rWjPfNctgi0v6DK+leMbzTfd
e05NfRe88DqyV1mJ07d4V8pbs3+Qig4za6e51X9fRI3FL3Aycml5jMO+WbtmIAmj+EJrU1VUC78m
mJiNNKqvS863ruKgk1XAyBts1RkzYBYDzpLPh1leetcf/yeqjnHmSMkJSfmZMszVMwnDsAe6zv6O
7oUoKz8NrismE+OYhbm5kB0ALWktpN0/tb6hf7Ja+0nq7TaVDmWvSwSTczIEX4ZVrui/hlx7kVD0
aVSTGm7sNI7osv2qLDrXvlyK7CHXM9GVI6K4DvXGU51L9aD2lkkH+HnxCT3g2LjIIw5JgZm57WLC
AQbDTFGIyPd4pGnSYpPguLHiA6v4hLcKfIT0XhLZVEKhbEZQs6kfI37ZM6bdhp+E+cVQYU72lYZz
QzTmhVkoBpn9a8nh+0z7QsshX8adw9FnuAZ08F7SulHIcjv2MSbcEMG9mW5+ojmMM99NQhC0BJtR
XUaqjjijUJ6TaSS1n/MeVmj3Xb9TBXDp/kTC44gnCsj1wHvVHfwTyb8/Kjuyu2K7+nh+kB4uHv0S
b7RBKs6E0n5fMGKgJgil7wkVenrgvuGRL7tEyofuV5gu7ss552WiWRDHxjjJOTiASxlMK4ubS+/U
RDY3l8yDcvAC4PaEkyAs2X78KiZQVlm3tYrBeHrZyqA3Jqh/T8pnQBGUXV56fpVkN7GXZY/ONcB9
tvhyTaY4XYmSh0KvwGCS/dwER6gRYto463djlCbcJSbLBfREOtVp9JTQ+6VcUF98SRzrBk6BpqVT
QToxGLgyhWfmTfcsfciq0r/dv7ieE8XeiJrx1118jiGY+ZNcgrcEoJRZO7QM7gZc9O1pr2dxfBh+
q52T3xyvVhbmlEayE8NCIF9QgAlS/7HUS6hgibhWg5b6SMy0t1LQAv/U565nBRyhHvndoTqfvgvm
dKbwn6L9DjAKmkWKmPV0ye1T2MFnTZncpIl3q2Nrj8pzQA0fPEsTEDQIdmcTBXfPhIXwNr97RjCx
fAGdh+uQIqCWS4v5iYBJmSHYB8J5p0EwYAz2YspjkRrFmGBx2DombcddDVE9b5gGnbRt+nrgtpf3
ZGEkhhmaFNP/Pm4d9sC/Micyfnu39ozBIgIrvrpPPb8X5X3Pvw8tr7dQ8YakC+h4EaeCLrWw8Q29
58AgRCR/qNKexKVAX9gYYhMAxVXNPLjkuOLR6S0Gu/cmZgJXQbSaWSa3ynjBRLvQ2mCrKfpwcU1F
86Bg8DGI0DlqpJk3yR9BPCdfKjw6NbLooyF2H4cOWhUMV0+QaRnjAUtPt8y1SBeQgv1AaEhui7dp
qxRQ2JHUqX0kpBy3o5gJ6xMd3NE3Md3nLXJ3oRC/+Zebv+DFto6L3/7Nph7D2D8JRZTcewzpSyy7
kJ9C7o+Uwp8KpqhAWfojzZYopqSHX9rx1cns5hfIFJKsBK+N4ZKpMblQW2LEhEQv0IwkQ1a4Lc0F
GuPtU0IIwsRZ7JPn2c8N8DybMxVuIqpoavzMzhsN3d6j0BJbo4bJyO6z0Ip0iDgtjKi7uOgufXl3
jBbZV1sHocpKjlKXKHrulAT5GhAaNM9DfxJ0Kjppp01spbempYU0HS6EpA1OZ/r77QfzT7rbSAeQ
QkrbkdawFZy8lc95DbmbrYCAB4vh2gpP92nSsDXQANepOXmb7g3o08NXjecIDCVyIulCJZAVO017
kHecPE1GMkgJOdnAhGB+5dhx88HtzJ39+YLGttihXDB2B+m3By3xAyzWJbQn7TwtrSoiRDaeONNI
3KxsIF64LX3nnQ3EwvoPEkg7VqNc7zvA2Z29dDowY2LkThFpp9QlAW1yw8AscMlbUYsNlm+URObl
xMDD3xfmYuxhmg4KpqcyqboKICGhvF8YhXF6svNSFx3FNQtHbzPXoNDiVOkUP9l2pyx8aV1OjiJl
0meZgW3si9JDbRfirdmi3Q37O78LCIhqnkHwarTE+aRutq3LpjU9IR7PkpFpJ//sTgGxP8Z1ePhL
S4tq38oZPZMPsRjrJh+Gx9xVKUU3C7JIVJkkk9ZDZjXWw7eE8bS4L/n1oHnEVdwG1mshvMreMW5U
vQ3eQcHMSTmNwH+RSLOf1AF4t4XjtTuBrUqQjkRYPWOHDmFSDYtxf2mtiBJK/7JLx0y4GNkfDI5P
bDmA8/OF4VjllH0ab/NXatYzhZlL/eolze3AwqT/DmPfhV964fPD1QWJfLimqLA5tNWwzE3NJER0
u/WF1YVxt+9sozVVDSeyFQVk/6RH3wIZGm/3oXquq/G3mohxutSqC/VKcudANmUdU24HjQXsK23O
hjkteg/2thNhU+oICt0wCdelljSsI3pqODDz5jWLI5Y8mzozGsW3rUFq47WvS3RH8Q27pGXDugl6
anHTuSCbCHkxnoAO24eAm7Gra37AO8weSrchLkXsvJyWKi6zT5+cI5mF0cvBQeA+NbNwfxcQMOzd
HDVZ3sYRjgwQ2soAzJHkqI3On31VB15XNL/W/jfNpIbw2bbYW6oIj5/sy76db+lpYZShSyShlZ8Y
rmbMEBsF5/oQnyN9A93zMy0EoezX7M5W3g92Kq5LQLRyw7ZWZZIRykBujP3Syfyuv7bW/TQ3SRaN
we8qXKHciUYl18g6gD/hqyDIi6GqcmF27ph8QuiNSZOFYTFEAnAihlqAwxxyIMJSH6W0GC8mpQNF
PYsxTj7lGz9wBkFdFBeMSdWXKXQCbIfwuPsZYFtk6hgBYDHfLxzYoXPBtHyCKG/MCCEpCDQaXB9z
nGH5KOz0OjmosB6Hgy/RTxeq9+7rVkayJlj0omY3zrqc2Erde9lOHCJyS1PUBpCbqSk22UO3Q/i5
SIraEJ3U0JrIcwybEDHF0SGYv8FDcxV5DzUM2DOPuOQzqnj3Zt2ctcYplrGP7DZMeduJPou62B6T
qM5WNKEMK9zjzleFrOZce5+F/pQ/FCnGUT/9Qlr6ByO6q8cXoAvbDeemGyJHSQ/Vw1Ht+2w5flNn
ruTv4q6Dg0uqabygptaI0MYvVOCpXg8SH3acaU48Iz0ZzxwEfHj/m94Y2oflImQlqKhJWrkOlkpZ
903ZlVRQ2xD6LJzAQX1QqPSf6RZvTO3u3EMrTSKr29T833XXSf5sNmGcmPHtTpn/ViVDY3ha5SWv
Z3bfofzTr+kWV83MyGHrIYtg75rH3/KLHd00hQUFIy8++uQBCOjnIW04/lvIA9X3EgXOS+fRGWxz
hr+cKuqfaJjz8CMvL+YmOdIniovGfvRmFuBsOm5q+EE8eLhmQ/haxsFb3wDv+r2l6cUYnUDz5Tak
UXHMp5w4aCne/750xG90WybFJ87ES0yC0WENWvBZ1/h8mNeW49nu8iX9gHnQW+U1w2y+8qWgodir
/n0Ozk/Uzd5NCrzo0qhR/rS3IQVFOGvP9b1bAayH2+qRKY720XLVyx0pbHrgkFJifFX3dZlpkgqr
Nd77EhDHw4Qvc/MzZ5xvXjQf64irV4zd0g50DG9PtrprHjvUXgonJVfEqjFwPdZRDyKrkg47Ol/b
iNQ0p5xdk8dWiJcBymrDBO5Pqerk9YSBz8ZMh1Xj1VCaSzyl+4r4/zzlL6myMeQ26XNu2bGlWEYw
cvtbzpRAN60J6ZIJQhp2oLqpUc5GG0FoXikzh9Lr74n7SdZAaBHnzqmvFuBU1W7HqB+95oW+v5wE
w+GB2h6sbieyQ8kKr3HI9lL+/oxz+2xZ4vKBPsTHqz7Rx5lzOlakI1HGYSDvhjwnq/DOmy8VHD2d
rntcS5fACpfIBasPjNgMMka5J0vrHn3ncX6kPkVUc5f5kP4eq4rEaqSGosQiIyJESz8ubDFNloen
AbPcgcvtzZcZ6axCNrZ3/0IqOM2RhYUaC5W2oC0hpbPwKrNwPXZ9OZRYTwg/9QikP4D8cN+mQuC3
E/aLiluj2wSKhm8pMz1AIdG2osjR34KraKjCfaCnyK8OSL3UDlqwAMGNnMqzpIiFs7dlldcWaPmm
CgDoK3bCSTcdOgyEofqWcisaiOCRj7/3b4vondcD+mERYH1+cc0WDBl4PIOKeyj/8A6ZJQ5yyhf+
4OdRVEVip8EhFjsCS9naVBdgMr7219mTnAA/SXD/Owpu01Bv0yftQzH892+jjnyM8UoFHP+vCRwF
GrVuN3jTrT9t0yNuFLt6VvPyN3GLDI3RgCun6t9z33Q2kNa7UIYtdRcsl1RY/i5RKglJVtbAwfOg
zX349Kn8urOnSMGspzxdwmMTNqw0Bit+OKUj7x6AOqxullcQ8DQJzJN0QgEILdhx7vXJNzzJ1NQO
0JJ+Ie6J2u/ezViSYtU9xHUQE3FrmiFW/PI7bnhAfCDvcgwaJxoLL+ATgl9UKV+LHkhPdpn6lU1B
OBssifjYaQA6+dbd7IzNLN/6L5SPLrdQHCQBCYQhaMXariPOLQgDCg+YH//TG34VJXRTlPiNjQxR
sWkiOQaO9ub/8Cla4z5dw7XID7Lz/g0aUSrMTWrQHbVEqChjrIGbYio4TsjsO9VWPwM6PnB1Z+Vs
puNq9xZ4p0UP9SFq2ADJewIx2j2oI+gtgPq6egi4JCMR7cffDfTA0EP63Ee6+fNkiuI3PzH56/j8
S+Xw+hhLeygZtjBhdDo+wGiCeveUSWihJsLachuf0jypQS0uITys921u9m1C63pQByGSXgLCUwaW
qu+n5LwgKDd7AIlR0xHpcsLWFZyJuFBXg4DXMzDGrSxZgkXyp5hPZcGh95E3D8/r9aRgzQe1Qn2N
vbYSpoB+vUDl8jK6gENn37YX34Q0CgwRp5EElE23TAK6WHAw1X+Mjcb6Hd6WOG9Plin2LCzPrytA
qPseruvDZgLsvj7h4wFqyrrfFSejzyxrJws1Hm2M60JVA7pwjyXZJCm3EaYUNPwkxBZOeo6B4Q+4
PZGdwYptqSQWI1liWxchB5bOZ+zoUaZHu6jEKcdTVDcBk2zEAXk23ZygOpnhRSG6S9KMBgnRUcXL
ni7IF+qFiqhRQTGNo0VgFk+1rqjvX5QKM73MmWfmXjjvV94J1t1VDDs8XWFOtSieyMrXf/vblIzg
obcxZ+Q70M7oPDM97B/K0diM5txxMg0R931Lri8wHRQ88oQ3RYYnd0W6VSEtjShqk3gDFsN2Ozgi
hX1AjlEiAStF0eECYnPObCMxnJIEmQEYYA8U5TCIEPr8KNNOPXVwwHfM4pZI/FG9ejCRP5nCRsq6
qWXhyTOoQDaKLhBw4esl+QVxB4b9wO2sTa9DnskhSG/CqTQWJBakL50fBq/g58gXArXDU1nOvAMP
wUayinpYW3/r+Ip1OxNb13vTC6XCX3AKg3tQqYQePSPxU0LY4fgBgtfNvy/UcZ42kRH0STroMXgn
ZZSqj1dfuzd0VfMHOzTsxqRqn17SsshIh9jxnPekGYeFow3+GL+ZE/46F+p3U7qlbDA/1kW1AojL
VtEP8p66xF8FOUu5zajxu6CdHvZ8c7ClAM/ZzqP1ckAc5CpKt6U2bkryGiEKUccot3yUpRzG40x4
BmMfvaycu2kC6XKE0o2iCfFY2/SNZgcuaXrxIdokceLQgqRgQqh/TLJu5YFxDKbpf3yQztTn9wiV
5JUmNuWnsyC382MkHUtbqY3ZkmEjQgkDvLuWcmo87nq7sZoLeBwKWJQiNgLGWOtMeKJr3Kgbzlyw
Pg6oqZ/69gaSOIqlMnTNYQ7VkP2fU0DiSZbSc/dAZEm2KwoA/GdHVoX9jZJcNkWMcGZWBKRag50X
HASyJfGE7uCheEIL0f3BcTEtvh6CHfbisNvDfBRGWqWjSIlO49l+qO1b/BDFFMt2VcG0VBiZT/so
+06zkecZbjggBWvi6UJ1B/i6C3PNvfCQmdHcZwVkQoLK6NnSJjysNWqa3YjiSIaVF0kfpSTEZetZ
tJ24S+XVYvNsukmtxXsJrLWfrIY9FXk31WhP0ZrZZvnWnj0AG5M70xVPiEKTG1rbr0zr7c82JRw+
UaJjJC1vxAG8OsMyvVTfVfjNtjrZHeCz7i/fP4Zwz8NryBnauga4BYtj1nGmRKWwPxtt3MXsAnJE
QnNRnr95rLsLOREcOvdAjBc0wy+OmyeGM/kFwyKB4HGTT9d65GY2ufCzAkKLZuUhFNLF6bjNjZpD
me1VIPFnPEjClDq2AMabzKfkb3MMYvnuFF3G+AvZ53HV3+9MOohJQWXE0jXbg7SiszlWs/MhP1xI
EbkrOphn9FoCUAklxVjF9St0Om5Vq0Zi5LMESrvzAhS5gEGG+MPn4SZM3882yR4zY0yvYAXTEIo7
mQ/aD/oV5vcv98fhKDLVclouH0G1mrJf2Dc1wi2Se3mBcDS2SHaAvzCnkVz84GeqHchgBihncHp7
CVWGPJrD3ydP8miuj4US4rKTnZlyZ4EJ9z0FG3HuLpVnwqjEadt3cqlOotoH8TmioW5sXW7GvETc
mMsGDAgFGZ4PBsI6lx8rua77t6HzD6Tkd8/cRfZLT7aGpK2LNVxKcPV37mSITfC+lgWh2ckexfDw
1yy4lGep6SgDRlctg2NzI8WXw9wUmBz8c6u80C+4T8EpYkxchk7fNptZePB4UL1PyweI0KBZCUWs
+meHZpOwI2dHeVb4tVAYZbSwkFrT5zBeH5zqmy2BZ1ASJGiCSGqyZWXWzbJuzujy3bEI5MZZGHTK
iPnS2bAeg+Fh3IjaySoWIGFE01cRa4HJfkQZi0bz0qbYayukibAVhGpxOZjrR0uXosOR4EVLF2YS
jQ4c42GiWSmAGfHt1ABxREMXZ65PegZhlrTrwTC6C5/lEwWEEH8SXM3eBJRknzFgLVxek/FspIyb
IvFZ7ZJsI9KFYPF8z0NS7v+VTf1R0RJ8f8tEv48FCDOaFSBxTN65pzGI7zMn95MjRjkYOrBzvaDa
I2FVDxp8RjOxwoqk0b7kbuOiBCvPYlKVTruWtvFA7f03EqI7i2q1gGgU3eljfs2gFbCYH59ymb4S
JXZTiBdYkNLSo6FTxMz4xc9GtHIMMjEqAzdqeS8gR8R7HEvnYvxakrpj7kTuRAIyh33qjGQgxhzO
jPPpDE7grbhu8ZKBB0DeXMLmRE+d6jjsYYszGvEq6n1hqfOHPKq4SNrkfikwfOKe58xEObGvzJP5
jpL9ov3luPztwOmkS5L5MgSpEVDHWxH+Vnkd7xb8YK++VDwx4pfwLEznCE8ZJYLai8qw1n5ce1pT
vKGLl2bogLoElATBV/X0snQYaxKYd0/mTMg3lOy+bICC16iLrLT5j/jKLhEDZ6JzOo0Mf0a2quRl
FQbSnqLW1RKcRchJgpyBFKNULPHdiH/YJayI2fPortY+ODRDuV2UuDaJE3u0HYESnwWzYbi/3YQ4
yPBGHU0ck5xHFSnlEqxz3Bg+lm/VzfN08AACNw3xlTN4h8dvYKkd6cJ8qXAwaV4ZPRvksYyACb0W
4pt4ZSsOmTfGAt9vYJUnfDnarx5MMzypq//KlkCi0qXcHIpIAV3MDzgVTALeTn64bph1hqrDAHMX
6ySo7OGXLsBVljlUtwj/etrtTqEkLWR4R95k+yNJS36kFUR8thqm7+6Wn7tkX+3A5zgGykZAHCKs
Q65KYR3AI5C++xTre1kxp6ZTweaVORSOwni9dtx7GzukoHiccI68cDHSrlJtls96RgeAqXnaB0mJ
BdFndJe4JrSLE0jkiYBnSzVL57awiAJJVUieE60NU+WFxbBx9ZZKcKLlcRVddZlZBjovGBLuVNhc
+EsKbDjZHQHhIFMpl/CkQgoWc9jQaZBLPB0gjFP5yXq6+FsjFhJSZC/djFhdDNC00Hocehfq0cNX
KmGm3tIupNDgQ76mvcwzmdB3Vsu1PqObUMnbJJMuCOMwoy8mPdFhLVWb0J2b1hzSeI1wnXHv/Oyl
rcMWQaIV24XZeaEPhcnzpqNOZ13Kd3jqNy22bpWYisToMNOSVApey0quYd6g9T875xkrisWl9gfI
DZkFOaLiu1aJeh6jPvdR2J9PfKk8Tx/xCYxGCf9Wj3L7zlaNNUnSjc+5rdGNOEND6+mvk496gERD
KF64fp6DVt+6Q2WfRM6w2Ducogw5rh65VwqtlVZ64+7VqxIr0wk3UfJ1wzIi8QAj9W1WF6hhENRL
MZ8RcxIJVaxRzu4HEW5IjaOt10D5VkuklzweEsn7mtHSFcmBAPlVBrxpWjox3gRmn0mH1Dk76AMv
yofUqCWfHDAP2+E9mtIhBwYvnjhxz8DXQCPhDWFf48fhvcvNMRXfD57q+rt0+ePGxKkfqDw9vcTO
9ucGgNmaNiThqGA27OOHJMLJPOIbwjoEQGVYBfqrlDP9vcYubZiZQLv/Ck4thrjjyqX+k0TiUnca
opVS4krhHPjc2nbopv6Lg8uIO4TI/cyFZxi8eXF1diZEfJ5zo7S3XOs/pwiVpXvL9ojFDJ0C65j+
N72c6HuD2mzC/G+8+gKn2jZEQettZztQUmtmNC0ZedcVxEx3u4xMdGk052CNXVy9VMGdmy9MGOMd
2wYhudpzBCB/MAwJE0uOrpq13EKx06SRAKV4Cc/BREd/xnoNiyO+btIWE6ZN7VIf0wjdZCuchTp1
FJpZrvbH9ADu7dHBCXszTUJZcmVR1RFHWOFUxcvlv8qMKpB8KSBo2qTY/EW6YPYxWzeiPV96a2oj
/AxaAjW+uTTcewI8ZvO8dZ2P7I/0JDsyVCeNNtb4BV5ddTk4nvIos/TgLlGPHnRekSl/F5dUaeW3
dZdjaGfFgyG6vmTq7K3hmvZN46V/Kr+LmVHxCL/saPxqT5YoDK/XQ9HPKmw9d04lJUd6sOHDiQUf
1Mg0m7/1qzIj2rARfwfaaoAPQqltAMXMFKa8U8MKkWBLcYjRDJAXPq668ylt5tVs2BIQFx7ntIC2
zJBoiWu1NEgWfAXCwZYCwCYm/ocde1XEjswY2JlDN6BTMoUrQhLrknj7sHNIv8LPX7oOCwheoGHx
BWZ3sCWiBfpNZ+ds83s7sZRSx3UOaSwt1VhUB/E4J7zZp7is2L2zQJlaWgmY/rSoyTDCR9aHNNUy
cC8Pw4cYuWH6vflpvR/Hp5pxEtAdLRKcctJfBfEfCtUH53C6ceCEcKGE8eiUMxWG+hDhhDr82RsW
0ErqBFZwGEuYjePzBK5x0OhfNLIP+2RXYQL9nF6+nZgv4xaBtP7OAuN/NQk23ZOwqyIrtkcvzevB
cQL6n+W/CJ/rqUbaamEe0THuvgLGRTQ9bmxmzXIWBqB8WPeLUr5TAssxDlJ7zcdoUJRjvTm9j2QF
W+lAinT3CFzmKxb8dOKDsq/N8YQWNZsB2NtNYhgn75GQ7L+HPhMvTmRaGLuatTck8Mzb/EQRQke8
LcI36O2NUBjfdCPTzDiG0icxHtrAw86S4daepBFIdvdWea14bRfnLBUep7lmiJCLDzzpc3b5h/Fl
miBITGhXwA8zuoNgnMb70n3iW5aELfrL3w8Q2nA6u7zejzhAmO2XgzEL6UDeWMdQfMgHCjN8BG5d
WP5XP5LVqcbp4bQduC19whVZZ9/7klmIV9CJ0FP5DT3+2lKUMUCgLJSMj23hmR18jCyd/DTFyCT9
zQ0xPIWI1c6ZDK6jm/M9F2onUYgBc6HpXMToi9Brylz/esSpO8Kim0St1dgyM+0Ha6Vy1zaeTYy9
OwYuT7DVn2MvYh6gy5SeQyFwW9T9RYmdXd8SZvQoTaSQP30PTGqQWS3b9BknnxS6V28ABnOvVMx9
1hy83kxj1YsZjdDsPieTNd9JrBXQ8Wqcfj02DEnuro3h42kFxqWVQqdrLbSpZk0Ivv4f/A+MYl8+
a3q8kUnDBBUV8AseItGeRD2PPoDy32s4dBc7MjAeZozEHfVlF/hLmH2p/TU3KIy3TZEZ2qUVkpRi
plRXls9b9ENwT3+YoQyJgXRjv7sUeR3ZcDYiQacPwAkjh0Ylxq1VZI1UXkVyT1AjnlgaJ3YEyhwe
I/L7hHPFyI3Bb9n5DNj7UmyKIRM5Q0AvNuiVzS85CPgiFbLxrudjrvCDe/FBV3+mMLo1dxMBDzTE
ZB1JJ67Y4/HG8zmDDwSSnQCPzzMmiCqubjweHcrNgirbFPuZeBy3OzfHfo6BW4k8MEZjtv4jDrgC
McRdbCoHMxqnLtxE5vi5WgxukjmcU1TeAeXlkinUqDrkslubCV/mda1Z6RcbY++FWTd0vFTuBMlM
5T2ceCKK2StaK11oDDbEJs0sNRjRWik5cmpMALKfO0wE1CjGXwC1oaCpVzF0CHLkwjAOOKxTF+s/
0E71U3MxfxuQt0BekXWmufLCeko26oyiqiSjrVS93EBTJ7IusYhPYvWiOhzAbLTuV/oEk98SMv6F
2KtZFVJiIBOEun8K9AwWBXoMJ99L7cBMSm0k6gGKef5a+uGmLrZGXPAleNuqjDNTCg0Ams6Cx2fp
QD2YTY/h2stzkskjrcaDOxVH8uKoSRnA/M8oisN8+lT+gONOt3N4MgMes4hSfWZf8AbEJxugc5gC
ZWqLY+7JjxQjn8xwscsyqYYNSfQPyPV04hPcdHK6R+XY40XFtR7KA8Mu9I+tJVicxMcnX2Qkl38g
5/7ueOnGfIJ59cs16Y9wN0hffNiuFt82ZKtJvUJEOiU/molRl4Ur1wBp9idBOpBaSTzIzHQh3Ypb
96bdFjgfoGIhKt9yP7kXLZ5YVf9IcIcCKR6LPUO1cbN5F88wrRKbKvwnJd55077h/qX5N+vt+riy
qE9ecMie8Tmf3RiLX7n7pgAxcR67R1BIQT40yAeuu090UiBlbYIqGEIx4cTfK7gGYyBRCKJYZhVk
G/fSF2toCSvSWf6/Jr7kPBeZgj2U2frA7PPC+lRRnwHPEoQTG/3rNS/WVT66PDRwB/Tp89OZtnEV
6G8EhfLVOr6+kR4aJ+2mpjL4aLOIh20ihjbWyM4H97exsQ28PTGqu6VZXYSQ4frTyc45bNWeBO5m
YxKbjhumsLDZDLhRNNPRZ6me8hOOIcimf4lNV85xYYzH+Tnrjl37tcq23ztapO2UGMUg+xtbLp15
sovozR4QWVtK2bFkMnOfnWXkUaiCdNn6iqfG/1EYIrKuuZOV5lbgp/ZsRog2MP285U56BCs0G+9c
gLmtFc6zc+U/ALpxEdQl4JcJPpMDL8iTBGAu9PIBwX9ukI6UuZvu+816NpTwKCd9cpmHxJa3E8a4
sP98L8MckUuq3qxqKHwlP5NhXWgJSISJFyWIpbrsnScSW5zZ47Eq97YeyPNSkaCE9tjCOlnCMhU4
oy0RLEo77rrlJDlWum91cagXNp/30L8CXB7EFlhVTXeXu1I0DkchGMFqY0agJrgCEGznb7RyEDKf
8ydmzIv7Mffsyn6dVx1/BLG8+8emxyty4IMuK2VrNcUAvDZMk2oIXyDUpM9tpqr+OE2quUFwrFrF
OUmn/Fa/IRDCkES9KHbbrvYLl6s8d0VMuBHWAJ4fhscx3f4eeBESAQG3V3VIF4mGG4ZjTH7JW/xh
m1PsNM3JW3XwqX/cHeEILbBVeppp5tyzISLfpgkxkdDzTEt4SMTGi893tWHWwFXHsTMkIf79t+dh
gSdv8N+zDLq6y1hbXZWxiZ1yrf9Y22bPP3V0iRvPtFr1Qdb7d8Ywhm6VVyXcZgONhpp2t0Qri3Gi
YUR5GodzDvlK2Q3Wq1gGL/t0gNzEDBHCWFZdIdil6oyc3N+9291w8BvfYC+qhmdoJSX/nJJZOEpE
zrexQDRz26j4UkcwBiyxcjrP2Bp7Lye7/HOKlnEMUZPdu2tyftZic4Vb+2n/2NDzTp6S1NOn7z9v
z1VEvZCnnz0tlJtu+PLXzZdyZH9PlCkm0i+mnzmFGv3eY9dTDROQu8fX+DJIEUKsLjSvkEPAjDat
gox+J1XD4s0+megjIeHtvoZTncPqX2B5UtmdvA4yjff+GXreSk9dJ8BVZ9Szh/8vbuwBILrAvNHz
LvRQzOWqgLFJg9g/unvPrU7cXvUUt/2D8jy48y0pI+j+pN3gq385L6aziyjaKUeKqcopee8+gA/M
x6lUs13Ao6lY0HP0uyyIro5O0iLc6GN00mmUqvzNpfIyJksWAhMk48FI7gVja251jOMF1JMeNA5C
sOn5qWGtlkGTzuVjQKNZVHNHQA+nBtySFkJzAA0uOt56Pz5yMt6NqM+2QevpI/OyDo2+7uxhqkbM
NB2e9pXLpqRXIRorazd0coOkP+9cIBWc5dLoMaZSrBwcTxnIsWzwerqpAoYTSftqDUFcbyjaBt8Q
0XYRRVaTeT8YaL5LqijXe0Vvk832f3q47/HTtCToe6JCW1N/sW+mLRDGZM+nLKgxmaaeLR68XSm/
2e6CoJIrQufq545O9itmjTn3MLyMEdeIxDOKQvRKWTFv4Aib2TtNOKACSWZpE7429XKp46DrfFtF
niMEH0bMIuBoDntHWFRJBj8Z89KJrfJrNfeZedrPdkc49YwSU9JJ+e9Rp14Nj4c5vunoSdrWecPM
aaQoPWN6OKk4KG6KYKunyrYUg5RfCHQF4jY8dFCKjdwnAquUVtd1wKKAsay8mD55yv+i6Lm2IsWr
4i3/sI8S0+LXSkC7l0giM4aHVymPm7Gcs5C2kcTt2kMLpN2L1++ImZf6KZ7SUDuHJYEdD00CgiQE
cc1/KY+qchIqotOhnLHkSQQpF76sU4K2dSvSNZidXz2AwBIrbtLpMN4vN2gPHBiUdtq2r7L7zEEg
wcCI8caruXErJt9TYKSGpxoGUEm14AoZE8/y6VkEhcOw1NXFmgjdZvBMB0lBHJ5qJ6U3Pfw5HqyZ
YYtj0C2RJIIl9giy+cINPy/R4paavzwydYOTBiuPSVteN1vALN0uHDUSdAq2Kb+2f1ws/IWhx7s3
gsTsWxaiZ/7dXDoWt1a4aq48E7n5qaiPOHwxWx/lSpMjZsIUiqBCOFlJiSWKKuE4QRttPft5u42V
ULg/ZlWJbvc7RakP3t2HQ/97j/PGitBxppB4RfqtWkx86A3v2NFh/+PX+g0liw1Be9w2zQeCXI6k
3ea9U5B64zmoi/MIhcGES3AhB9SDb4wG8RU504LUvkNyJToTPl6PoNOnro/o10TuUXXmhe+W7qfu
ggiKmurCY/FAwBHOVAlYHv7JhbqfP4i/icMBBfTTw0YnChjj+A5oRRyfqa+i4knxTjPX87MhrKXE
GuS3cK+lOywNHi9Qr27c3Y8yFgokFMAlJGCfk0POdmTE1TTYxWfXt1pinp5km+N6F5pgF0Xo4e1a
zX6JEZFJpf4c69nc0UO/gaZ8TrFNP4Um0Q+CCH5qHFI/TlvBGtfSd4cllOd1UV9GLAiEIE7ALd7Q
XePlnlB6KHiugVtRA10WJSb6A2z/KLOYR7g/dmpX/hMGJPJznqB60WQW4OT4+BehLAxh/kbG5eLr
rH69IqCqJdNHOFIdE1pYUp+QvxKsy8eiY3DlYO8mPuvWPhvwfczTBzz739HuECjVWDLfTP5LHLRH
FRDlmJPcDfSuXk7afbLaflGKgr1lEXaoH4eBs24sTCwjHWiDdcqht10r+SWkCbq0D0OzWGc0aZJm
qcCc3V/mpRBHCKIETJRbAb8dhTaMyUoCia2Hwr8Kam5E8yU8mnbmrfucjaxD6Q4xdSYh21GHBKz7
e8sqAN9C9XnW1RbUl8lvzidOcFPngO0FchD3xR7MkAyw5dyG1xM9Y/iPbfWVfKKM35TcP+3Ooa48
eFg6ikd3ihgQ0g7kMk44nn/VXysfCOeYK2zWr6U3FlEMfZByufYYRSNHKrOF0pcdY2zvTIHNJGCZ
+FcGH1/Q971CCbsU9OnbFCPaKvLHazywBQKoNv3sF2O/xH6zDoK3KpB1jjbz9/wNzMWsUH9H4jv2
nUTUJXhIBe206Ra4D39Z5fDAlqgSGssL5rllJWa1V2CLCSb6LSDHW2//DtSkQBFVNggkGU1gneZb
1rVTooteoym6oqHulnGw+PT7ypMxvmaEW86QBVdkioMqdHmpDoTi8MWJrSpw8UFc9dbIJ2kRMUdp
THK2p/PytxYxdLQmHYF2AyM/8qQwZyTSq8v+r2j+DTsu8SMnp63NzBNZc7a71rgwVoNyJr3RpaG0
EN0tqD1NNBgSv+e8rDSCYIpeu33TqdIJhl+u92icTErFGraRQ9n5s0t1Wwf+lVVdHAUli0N0mUv+
wv5kskWz02+ESPTuEub72P0kmKQUVily61auguvIS7ZayCfUAkf5K2mKNg7Eqr6UG3N+rERmyY4M
IV5kiObm/ip7PwmkxlSSlW6+NS1HxG5jYjem2myT0NrGkMKJH6OHZil0TysaAH8H7Lc2VRRliKS0
MdddbXunVrKtyHRWIiGtGDvCWJrskCMJf9yevyaPWPXAFWAQkHYkj+71wZsi1X/injuS1OyMaNmb
3CdyDR8BJr4xe/Z26TRudWDGfq1kcHQE9pUuyzmHb+bQ0Cka9YUBcv95FPVAXZHgix5cX2D7uYa1
Utkuc2m6wdFdYuTi58fi4bYv2tY3BM54y0kkBS73Y6s8H62mRVeFl40ck3T0+bahUOBQKANn8FhP
crIda2eCNMmmJw/sSjgSYGKbEBPCegAPpcRdo70gH6fGTWXo9PvyDxQ3DCL1hLK6oZ8vPeB639bf
hZskxYETvQE97f2zQtUviMIB7ZeLWNgeXKVEbhNRRiR5A1zJKjNbZDnEZH2RcYiEdbWf4/U0xHKE
vCW8f/RbDMfVW2NE2212ciAqNLlXictlySGncQCMMK8YC01Ko57mLrLAe4XoSzcNe5ZvwvwqCyHW
dWYdkFTV5stj/sO9Oh6nYnxAifipWFtL/17sAZ+r+kAzeH6+5DkUToTplBMpqwrKerDCoF5FL8Qn
sj4lIEBgjNehZC6ZDkfl1dfZ1kBXOwRjZU9V0ZriNi8phjyPoaeAjLt8yJCYdpUK+rdIh+X/IYWQ
jV/Re60ZBhQzDwkelTFIZiaALpgYOo96EeeeBZPPBXqy0+DB4BZRk0iqIaLyYY3sFCsH2nnJS2nq
pMZCyf+02iia1dASbkKfTOq1+k3Y2dfjrGqeZINr6AGMG9qg9q8/P5vCdr+hgrt9upD4+fo9WFeB
KTCg6uDnxT4SwAbsgF7nZK6g4Dnr2HfOBvmTQ7bDbHCOTJUJaGOrW0a2mU92CeUP77/aWZGCqIsx
BVJSikWmsp0SEyA7G1Z5ZHsDvZvg9zS/ef20jn5001oEl+cJGHf8Zf1WzTWhRNCZZ/FdhMdpPUSm
KV3ouZOonKkx4C0BKbL6Kxjo0TALNeCbWdXwrRoreW3erGMdzzw29IMXt8k327YoPy9lNbfygwWi
bdIhEoejwBHBNlL0k9Cmz7AAvIasb+vaGY0Pc+XGRSy1OApLGgZXSsFmFD/oOAARlqxcoOA/m9Dv
cSrJwYJM4Xxji/JmCOmrnxROGn3R5cWabQmtYbGEp2Cqq+7bt9BfF3uvoU7KKveGu/Vtjsr0boVh
TCASPJlJepV4fFSuB3wwLLM3pbFmDIBgS0Mp6X3Z0Ohagg4hNKzXKkKs3E/a+1K6UYevElR5s2hx
yqv9nBkbFTafE53NP81d5yO9oxl2g0SDyxyVaCfRSFLt+QZA8zT9VOsG8q7id6A+fG3+59NzB8aA
mLA8Zef4gMymr8TzAbqh8EDh3KFIztpO/Mfy+3nGyy+xLO5TPvt6tT5QWkWiQKTYZvQQ1xRo4n8E
Lm6Yq90pFsO2UrfsYJFfqJBf5KtwGO7OEnwDYVXlw8o1dMkgJX+/9oggo5SVRUe/I95vZwymcW6V
Ej0iCrxdId6wQ18i7/5L313BX08ysPLQc39ZwRqJ7yTrnYmGE4PUHnsk7mV6W7mIVM76M2nVUx/e
jqQwoc/KOQ+yQKMtqnyfx1orLQYUqbCAwl6W2BqTeSvxIxd1KrJYhSc2UNZ3mU5kk/9aW/QmDTp7
EcYpN/dtti4VPWzBTqLCYn3b0WN0GAJqqIGCPJag12UIYyBvMxA9KFlbmhja+cSMtXAooJDDa+kl
cuckFYf+/cEy0/F8CVxHZlDPNpI9uyCY4N+6+eo+PRoQrnIPkmVINLKHA2NrvO20D5JjGA2BbDZr
Vq9GTExWsoxzAcR7cVK4hTCFeDgQeCLyC5lJnYwkeohF+koUBQPBFPJZVrWuw1gKRZakz926znQb
wSj56v4XbetXvshA2Wc0MnuI8BNE9NZCm6CUW7q+4CfPJ8uaUl2nFI5J+f5kVKo592QDVRtJXEuy
nwAY/ZB1OK39DoGT9lYfEummIdLwFdD+YbskECPbQc7dSxVzGuk/GuKb1cG0WosYDY2FMgiSFRoQ
jnRBipxCIb79+nWqAZKzgfj9zzO+ysNLuurqNtim3JCDbKrh8bB76hB+xaCvzKBvWta/GlgaXdcN
qcoaLmCsPLhubCj84vRkmI2Cwz5AC3ehcsnUCDUT+d5Gyk/hHUWTn+5An/TLZXjuCuTRA0m9Cd5v
D1aQM4mJ93LkFLGhwYFlEonUgar1Ag0CCIA5jk9rbCcYyS8AiGxsIhHl7PRsRoy5LCBAe1m9g/II
RXSnKfVaEqzuAUEQRpd3LVX88iDmWoPdTmGsYk6CgvZer6cYJdS2LvHElGkcIErtr08lDFWiULx6
jTUxJLbXIAqoYgvau4BjRZA+/q+H+bvaqxRmyG/ts6ap64tHIZBMgblCc70s2hsraKTXi4p1ZK2q
SGmavj3Vr6Rfg+0g3LG3qsm62Z6zuchpjHOAilLB6XoniI/LhiFtS9c0eIy1YYmsm+NFQsiw6i9f
Z5cSbWDw3KIBJ0Ejw9G2Lli1CeVyHu9a6eYcpIa37WZmQzj3kHfBuOi4BIsOF8lAaezdRLG8BLjG
bkIlNZRfIDrOGStFbIVtNDmivLoQLl8djwNxoBbvAp1XYHcIrPGUPSXUWCpiqUZwXth3uIf9W3Kl
QSTGOaJG4AqPHFOX43MMDvxASZQni2xzNl2YiH89CDEgyOgx/bQOuBSlaVg200n7pobnk8FGdbi4
FedMf8Ua19Rjk04uQov7XgLyTUWGkxSpoaFvQ31zP+ViXv8ylbHgcZ+xleGhMNuQ9jskHup7lxXs
a6u7JkGQsCtWrXrEe9TaIDKTfjkC57JGqDuc5WbBRSMclwuUV4f3lPPH+iezoUy28/N2UxEm29Sh
TtTv8fv8UdJ7NEp6PZEAvSSo2Ee05cUQjWTf3Q1mS+qUjgSs1MOv/LU41XnSRZvCuT/ntlqDnJun
+x+AkDJoox/C43rIkALUUvTBvpl5MVoX3wd4C38E5D6bnQQdlek0mUUvT85hMq9601J0dOUqVka7
mNLlU3CKrRrwOF9LyUhfgju7DNoezPq54bstyOPaP/+NSRlPZW0dKvmxNhmTVLIfZdODzT0j4X/2
neiHvp3v/mD4+Nps8Vcot1S6POinkb8i5uhCAP3KPY7NuDjs4/7IIM/+qjhBg5JKHSF76+XSazLc
KE57OUDn980sIx65v2eWXYoCxmnwawIJSRRCadCIP2VhR2XB7tT68NM3WUedlh8cDvaJEpWm9Lda
qg2t9aTcxCrIoyOyfLMChHzIFM1/3efOsU/sDk5/5SJkuIkdpQ71sehM2Uth8F8HIWCWCqYQT07d
ZyFMnLZfvLcan+5uWhkOPhzXIbV24HttUiEIo1HLGmc0o/cN36JsEIZD00vjA7XQaa9iXfIV2IlS
nmu7A1pc80suAKXN7tgswSBxESjQlBoKn1URG8ng1QZh/KnVQB574/4zMkTSepTA1+AzbFoZ9u+9
oZn7/5cndzLo9rhf5dfKww79Lz4JdI7I2Osusp8Id8jgMTcam2IOr05CEAc6Do4+gXoIPABqRVS5
UKp15Z6gD6W1mMJCSi+InM2lvpu5/n9QEcrzraS1pT/PJfES/0NI9PY+ZkGp4iYCdQIWvAG/M+Dp
oIwHNfz20g+EBFqZRw8SLJdgpIkR6uPNZPNMxgs1GDC8bFF6STnCQRzw+CbZxngs2GrC+pzpQwFp
+P0+t8HXN9/v9WL5aGsPc/93IlQ5sptDXjD+QORrBnerayh160v5eIQPY5U8XRQAP3gu/4r4kbnf
vKc4cZBQfzMdblMCEW1v+K5eU8VDpE+T4aChcBGJEV6xsREJ+CBPVbzQhdb5S3z82LtuYJuVc/YR
QnoAgLKmXhcnC4NZv40O3NuBb9kpVksbcP5KyO23jwmT7PhAtz512efrt8JDxI2oUq00TgD3W4xc
3ncHaGh92yLXw2r1dq9kPp78vKa9ufEMhiLRKGFwWhXoCgrJOYUe/UmmFsSpc0lZ+2FZ1CqXyBq9
7Pb6k3jN8VOdv2hA3ZFU2pEGelSTgQspKWtc/gn5S9jEjpbbHOeOp8jvolZLY1PeevMmi6IxSrMv
fOdrwaOCeQpcCWmnaxt4DBOIUPNxcILg8jwoKKazc1yp+l2PrjEszufVhmnMGKLwsAgZCjOEgIS3
gXN+n+3W7DRDR90zaPR760nkuLEXW5f4zYIIdM+845BuMoih9c77D83I5hBzAzGZn4cSeOutVFJJ
BZHP9qljcslJT9I9Pw1KN2oEqXXFI7jk6WgeLuHGtJumxv7ZZ/p1RJ3yLSuyDhvacuOs4UzA1/nJ
WNO4q6dtxhYqzBZkm64Og5WCTqv32YmK7vVapWic2AytanLPMagWECZRpZ+VRVLJIJUagXP5zmzm
LRi0evdnOR8rC0mJx/AzHFIZrkdBjh5QXdg+niAGEX54zJpn/ztJB2HXKu8LnQ++mXvUStqUNcXH
GxMC0gCWBZAicsuuefi+rIqmexLdpm+cTll0pElUu2ONcuARmkzU6bzTlCdCoIL8nXftUQd5UiBs
SPfyA3ZylbmufGYaz7h9lqfI09MySsiXf/fMO8cAr21LoiQvqKW54W5vsRFD2cf3ttDjSfVnwHls
Mcydy+Wq6n2P2Fs2jXjvUE12+0Zjp2QJ4BFAa5VfITPJ5YXFUN5CaRqF7lAxZhFlkfARONM4B7FI
Lvj/w55abXYNQkDQybQqzel2qgQRiguJW319NiidUVDf92oqfmlBwrgUpHQaDUFXqjqNXB/J6EVU
GDO8xZo1mAwGXG/2vXNldnD8U5juuCqHjhqXeKoEqznAsxDOKfYU0S/0YfGfMzM4tPNrhEnLW7Yb
HOMlMq3YPGDoUI2WzZw22sqU7Cb0UQqMFD9Rb4HK1HXqiFeR2fiROUAh8HM1rg3D4tCrD4EixR5n
9iPudEILPr/zP4ovIYqFUpJlsoToRhAqM+3pZaTEYgWwRsUxVkhj6VH2jdTFolIuebYbtxDXhXfP
EyJEVbnha7+XlhXDTWxQWiIYv0/doA/PdZ/bRs1NI4/Owp+Qw8QoW1D7oh17ewqx8bKB0Ih4jsuC
DsBAdBmqQ7d85B0xvyzRg1jcFfr8I+fJVCI3eJYxcBL6plT0o/w7ZnaRv2Uc7vAfc0LRTZEgvAP+
xIeqE+z/y62aLQ+Kp94aJmFCNYSCaUEcBGVXRiKOogW/US8HcmXJHQv0WBHG46ZHaMxS75SIo5fH
woo58hUF0lNLh2QeqbSiX90Fn4jMTkQY3rGCkcIKX9V0QlYMK78KwSK99JBOyjrnhND822w7IPN7
Rmcra3HHMgSf7QG42ijUkgmdRa4TnG/9j6kggm0/PXp8qz/2vYIZRrAjFa2kSsA6xkZKQcgpJNLD
M4agga+DclIMJzw8rV/Zp4nOak7szCGyMZkkfs4gRWqmHM+Pb5eFxt8jm4X3Z1ITRgltJ6wdLGDn
mgh0EWhHZk/+cfYd82hUSpzU/Is+52eV/f7BrIDYReNtYaoCcLEjTNwRzJf9sVmp9dNLHdaLHW5/
4GOTAA2DhZKuLQnsKCKM+XKntjzERvIvGJ2KGmk8de+lJTgm1r7mN5IIfeVAn3zpvrMhrINMn+kH
fTXy89R8DkzR+QhlUNO3+RIrAU/O1eNWFkCftUdBuYcHmD8R6AV6VAgJh/EdKhzb3O/vWy4cal4t
7e1v2vNQ6Mv94oZIWQanwuTIpekQgU6oNBJVi2bhtNwJ8UnApbgV36aUND44WZsv1806l9V3M9i0
8r2Py5RcKlGHVcNS8rHynxBA471n6SVz04P6QYpj9CTm+8hJWqqsQpwX5ztKQpBkR/0wrbeqJbke
vWG7A+GavDDdhmyvmo+6r3HOPvmbgSLSIhAvcqCX7h6JA+rd3J6b1iKujxpawqRJgi/wygem8/xt
DNMhXUqHF9/XnJ3X/I/s0a4C8sVz/El9ed4Wu+HFJ+W6C23Zp+jkyImFcBtGYBJJT6OJJty0AliZ
NA7lNO+BatMCDoLbkztK6C1BBtv8ei/CKBACb+2nRgdqInlyiTVxMQTlU0i21YP7HVFQ+MnkpbVV
znJMzYx7DXfADQeaate5G7BhgNnIsk082nWQTIR1DzlrWNzEqe11qs3EB9n9kN9IWbEIxf/AjNf+
Ilx9Ak2b6s3erMYDQB0fMCi3v77xJDztzC2HQdXbGUQ3WAta82buAgiaLt4/t+vG7Qs6zm3dNWZa
HxYVQXb5MIUxUjAUd/wsE3b95PFBBhLgu+RIGtFfvjhjt05NvDXXnMZCv5MRfTgiGwr62oNY3Z8u
C49zvzD+6R+U6YXfoH5wtlMbmoCFTNM/ZC6yVMc/qWSkEpkvv0D5f6bcy5olH9/nyjmg3YZaJ5YJ
zEcHVjYbRGpIbqwUUKgjL9oeBsLxJIEf2/MZCuGGOQ/9YlOyHL38lQymxIJwfiLFBv/zHoQ8VMr2
cJytQ5pI4FrWLSvHdb9Natp/LDgZAZIUH84l/vwgg4K1+l3fbKg2fjjuQS9h3NLNpo+Yy5UuOcCq
yk7K9wgDkWzYlNvJ5iwtDyCaiW4NSe71cOORuKFuWnCwlblvwPIXOXBUBh06fVL3j+tGieR4HchM
4fIs6ja7p7a6BbU9iyEKpKiqA76q9QgvyJ4dYAzklP+jQUuZ66V+qkT6UxKoARYuHdu4dRwsSCUO
0AXChN+NfwLKZFqPRv4dnzKdEo4cSwIrHltOPXOHEDjZpVhuNaByuGwpFF19AD5sR7MRAKyubqRi
uuHbGHB7IGnicWt/5ITxv4LY4jDzBWenM4vb7gEHhRw+3mOxbb5cZUdSc7vo2wJoE+GDr4a7UIb7
bFPFZBo0jMNYLxiaf3aX12edC7TPm7DzIBKDdGYbcMsKn6PYIUTiu+9KbgAFK3wIykEz3qa90FGf
M6IqaqPZMzxD1eCyi0EFwFuvyI8Hnqi/dx53mJER4ATJHib+0s2m2W6/uCBisUfpZfPIjWiCMEiI
v7wg5oZ5KDOGFnMBIL1WekdXdU3avsWdhIGDydLUNqqznp2GMc+N3hxFuW1kLWX+3nUvdAD7oefK
3nS1VxWUhCIk2H4QzuPDq/ISNDrqtkIVTOficYLCtzqOIKYAInUp/9qTEF5y6NxXw5ew7cdf5/NM
KyUx0bbqcv86YNDs25ovXCn7ZyX7gqmNEPO/HldekNDehl63Al8oOQg7lqsfH6LFsl2fiBHfgHW1
pbHtqhv+Hg1xg2KUxSNrHhvLT2A/u3qFEUwwmygiNj0qZlDZ0hrY95hpoxTGJ4V5TpKmuTw3nXYo
FxMAzTsnw7GTikztVoh4RZfJP/CR3CjIMEGdG55s9tKakxOiBVTxlJxJhTV9mVhEQlIQ+AZ4148u
yuO5/aPhKrpDD/ACODJo2X1Uk8zGqoNt3QiNWQFckki9Ep5QbeRMGZZwUyNt/xSFls/olRcUNYE6
BRxaaITDgZB2v62Sxl2KJEEq7V+n4PU57B3nI177aHVL7OLDE1yMEQolV28BoAVRb2NAtT9f7LFv
YisjZF2q9FLiaVqe40Cf0Mbe5rv9sT0y9IXat4OLCHeT/6d7ftioc6qXFni/649ZSv0iIi/sBXd6
Btdqq/GBCbJ47ibKzZcwFEZFbo6A4btMmzf2qOotM+W8YjfTxK1ozB3KTzUtKSEEV2IXFIG1iK5n
YFO2PED2VhqD3W/lTCHBwHBDJBcr08ltKObUbv01TgGlgaoS0zqPs2V37x3VrB/41jawlc07aawu
Pl684ojkM+IzPf/6FZCZAVghy0fN7gz2kCcZOG1WgvrqL55cOuDMSJq8nSkBqRhlQRQYncuC+yDL
RrBjBh7STQOWz3jN+wwgKaxBm26SWcXm7cePr97gomXxdb5kFY81RYgW+qMcS/Lueaj86/+vn2ip
UYDcP8T3c8PQSRVEQyYQvHummxkTqhWSfkboeueJrLGc2qcO3gluFhs0GTbNDCXYZhtY7fuUiy4r
loKwIvXEb6YT/wywn/LpntAR7uy+kv8/KL/5xfYj7xr9jJ8bCKV9SG2u9n065Fb1SgwPdsz3ne5N
rU5JErT1i5azpTcyDDlmsa+9YsDZgH2AASdsOqUri4QPYpFZo+plitWDdkv8k9gJdFrIfk6BM1bE
wp0ijGCRqBZkMZYvpGBBp6JdVBySS2ekq7IRi0thL3rO9dMYbStObH15pr1/N9zn0lly6WXaRkIH
VE0Qp4hyoPYMEsA3q0FzRuCDY+F9gRY3Z3uyymbiZlIJNxPPFI8irqpWhIQb5S4RVFQfL1QRvqId
vMrZicM6ncPtaEF/dNZz6oqgSNYz7HYlpfk9afJWX6fx9WoYJiiBg2qIw29fM+qxlEErpZtW2Tlj
WjrIZ2nhkTLkFTW/fMl0a0s5oA/gWsHT5YiOhhpbHRRmNaxaLuoRmpFa+QM1ucB1HIJYqgKyFEb7
IcGu6SdoymM8dnFvNcWFUmzfgG57lQgMK9LApARXUrDRZJyTQbQAAzfcpTBcsbRcjnAyYiWc6JLr
5QuJboKux+AoYClR70TR8WiJY8j5Niufxb2sw3/Oprll5PwnofqEvMapp/MjIeunDYzvn2JUjdjV
lGJ2Ez+L2qL6CqKLmeTbUZ55LktmcjYVRjgWelBQiKRejASvwrwuGC+1/BvAYhdDBYhbD0wMOpEN
XciEEZd5mmzbXG5RwLhFzFNZHnA9aHnGhDH0xzpIvtnm2g7lSrSgKM9W2ijSzIgKBjgN+C3C5qag
dGLevd0hkkntW4CC8FMRwi5xmbP9DkgPAH929dbNpxULrB3x7ZaeqeLMspUUZ9rFY4c0NvFxjiLZ
JIsYTt6LJij0eUb6azZc7Q4pWUcfbyI7x3UqCPr4YFl/uBVOGlVswcG1YlSplGW5+X8OL7eWs/nf
Hfb80T+6+3zhfh5tOJyo8xLF8j6ZlNDLyCCbvw6pqlbGCtwL9KrZBeFHNzGs6/p7uk7XkZGPeydH
dQIdrOHAaOnFX0O1oMeKKIDMQKC4xnTBCNu2Jl/ENzxg2yx4HNvaDoPolGlywPKa3s4R7xGstbiQ
7ggowwduGTClmITTu0ZHbe8uTq/Wu7DPJxbYyZhcX6QdU+It05sANMf8XV5pbonmRwV4imNvUsOb
Omz9bQrFy3oXK1sMj3/ORWNc6tPGbsV+kv/lhoUgAjhppVTj8CyTr5SihN3RdM4YmUIEuyzr3Sz/
7TzwLg/JOt//EfFMKTI9q2DZrdNANK4KqFPYkh+j88p1SyR/sY1zH2EfMd2qM8U7TI2EznKxGZ5c
stwqcB8mjmJ8BefAxxh0a1yFQG1qiYhT7gXL4fE6U5TzwzgnrK0TbYZQt9Eb6LIMLTB6k4NbWeKi
xUm2Wyh4sDTrY0mXEoq7khnghJZeeM/9lGKVHJqvGlzsvwSWBA0Z3K79lmnT4ODb4sm44SRrVXqO
+hRi0w+xrJteDSch1WAzNjgffbwJEZvRUuomiKTjfMEiP2mZt/VMtSYQ0S1gOag99AA4a7M25zMY
i/MXeyaNB40WfKq4JWhBwKed6xtU21nA1Iw1Q4CTMtJmBr0JV82ZvMOVkuelPPHd6QPdFShY+XV7
uCwxYsobNMlwlT3NJZF7JzXX2Arxc4JG0Fe7WBvBKzFrJP/qMAa5WKLiDCrAplckD/HDGxOItbfF
lX9f97T5tIqQ0hD7LY+kIzkW8TFgRgo+U7t0xzVHj0yrZ6rIH1KtZMvwLJoVjRzAbKEK3m6FnHX1
y2wYS2k2Jqs+VkFK0Wo1Xv84MaZmHpAkUty3XWIvyVo0D2lDPRtVowC9L6KyYrPCXrqAkq/n1eUV
1P9PJB1loJAnUR3D9xGdOdY0xWBvBMNkgXd3Nd879h3KqeyJlSLWyi88YXA0ml3QwZHP2TWbBmPv
1WdjT0gkPDtLrUxhc8Qn13JcnAhNHRWbN8lEXI9n0pwZx2ZihATcBEnds4ne9i0wnPgBd9fhzJTd
zcrVllzTy6fqNN1EQ3kZ6cTl/hzuL8VJm1k2Fnqayb4Nv0byuN+wgXFLHD/E+sD4jIul0FQJYiEJ
e3NsGLRjfw0EeaXOViN7F2sQg6yf+L89ZQonuGs3sgLjBQc74119N4KQRyJL2arFKYeIvcKComJ+
3vBaceIcLGTRWF0nWos9vc+F8rdtCHQeEDrdEZg0I3D5xaZWuWXz3QRpFxIj8v5YHVgiHdwT1Tmw
+cedqxeAUSmZ8SVIFGK83v9q9vbkVSOdL9q0OX9Q3JFculB8j26hWIJHaUSRZ2eqOOOfrBQ4l2Tq
DZAHPTzLcW8tkCJZEkTpGhM/rKePMbbpmNi+B83fMmXoeH1o51WgdxxBfSjgActIJbt7r9EXYhm2
yOdxcgVBIKG29woo3TlzKESQq8IbPIj5sxT2QlhfI2NxQpWSqhVn828iqAwd85PZCD0v3IZBugi3
6d/FCUGd+TdHMH6vZjOwoyGyworevT0FvlYlfTjTXs1GHUA974xNGcuOfo3MtEFfPsV6W30HgtWW
0NkGCcb3+IHIZqUWKWX5wdk7K6OkNb5NJnUkKDwrgcy6ah+dGNaPG+639gfmtmrEt33UHUiL+9/e
2WQoLUc5BCwDGQmWlDCcj4055IHVN92TMusohavENOfpluv6R5NPdp/1LNGg/LMhLyushs26/RIh
g9AoONzoWUriOhmOEpJIr9ULGdnuva9hL4Zqx0m2XE86yo321MjJ2dgdxSk/t/OUGt6mSOCHXaC/
0foXrEX2zjkGdvpvKalD68qwc3fMrLYChQwhDLRiWVqZm64UXfWhXv3iSYhomJ5t5jNsHRd5hIgq
TRhnW70WIvbwd8uCaUIt0n1GSYxPG8TX0llkj2dZaaKBqpOCw13KoiG27SKyF6DqKCFZig5FsU5y
LCWokbw/HQoUfrGhm7pfpVktRt4R0V+o89a4fyLBcWcfDuTj8RBOAJPqj714A/eCrtaMd6uGdt5e
q39cCpAuKB8eZgtAl8NeyVLh3SQJCILeARnuzFLFg6D1XJAg8v7DmNvFV/bG5O7HloguxQ68StEY
SVIyYK9NVTa5BE6i4HI2PKnzl1HPimuXH9sVynUENlxa5lnK53xWwPB7g391ka/1HuxWt0+vrmw7
yMMLh+5BTLLJoXGlUTZH0n1wGWnJKZIiOOfCvTlJWNlIbIpxH1eUjPfohBp9NDv9QwxlmEvFrWMi
v3nGUnQuVgbBLgZSybQK8dSHWwt4VXL3YJvyAwacNxCTsJ6zasI60SIyP2DPwOe7po3N0Q11DCdU
4vjKdeqJj3J6z2IS2gBfwN+94y0uo9in8dPzKysC150sClNH4qBFWDoh03AOWMfHOxEFamIOt25W
zkX1e26emPgWhcdwO/+ia7stQbx73UJeQsg5UTuUlyH0kGusmnOTNq32VFhH8B6gqMmf2spsVlfL
B6Ra2RBn7ZEmdHMROzT+A6cgoCgijqTZpPLV9F8vOx9BniEZCMVe6JOLMsuVydDNXruUGaGTzFK5
CaST90uhIh3fra7RUapMSoli+hcwYXSgTqmS2poQ5UduO3cCNY8vsvFV/Fcd4oJIOOLTN4vWGiCP
1wluHsnTtNv642FEzYZAmNS1v8bfZfR0HBbiqvTrkC34bwPHhr1NWiTIBVL6+Ym1KM/XkBnLWjUO
2JxzmSSTiTdPQmN4LXRd/8O1AEyBztiySV1jcpAIJnwfUqSjvSOS/LZjwmpq+6Ti8TWjfy7abHrX
p/YJihJg9MamnOd/OG9KYcDb9E7/r5ZsdnxgHZUhRDjVoSoCiMw/WxK3IVGJ58I6QjvRVQS04AnF
NjA9kijgpszv5DygSfZMXAG/kOmq3rAZg67aHbFBGjwcZFCUMEbP3oYn/YnCjqlniMu5vPjaBqxk
arbAz3vmuPosuXJa06Vh6zPTOBQFStmmsSHtVQMPM/rU5y2NzuCFJpXvHvUW2f7m5m+yRzW01cgY
fXjnqyf8cdpmWQujafTqtw5HBsVePzqtJl5xZG/HWFKpELSDs+t1Z2r93+MkxH5mgpPgPLlE3OeJ
hINMEs0MmoUDMsBUMm42XeNZywNhwrL1ksFI1kkA3k92uFAV9di0A9UJ2+YJ8zX2xEpQnWrPpVXl
Onnbv2F83YHVO8TUAvxFXxPLq9grgHWV+xZ5stqmqgqH7hyyWy6UWkvrT/PfuJtXFjhPwdXD5GOg
tV7Kx2zlLVtz1+hqsMzaJK0ETlecdDc6YjQW2GizdM8zMjhTuuu7KwZk3YZPaEMYKo0opJHrUlKr
tdOc9iXkS8Bcs4w+M//QvjMgS1yJh3Ei6FdkKYIhrvKRi7GcwRfdiNOHvv3eoR7KnORm4DYrnoLc
AXwnODUymvOAQlg1QnvzXtYz2UKjbNnxJr0vFjgy8cUKY7yyDtm/Brhq/aSjUE3FtU+wCOBc12JH
DIwqwK+KaBxi+pjyV+XxfOu6OiIm0+sGmZUjLukWP6b1V+MrcWvSAZGr65+fjjOig6h81iUdY0dA
aoR2zAYbvjjwbnoOc0FN1Xyr17BeJB4q98w9Ku9zUCUlyPth9cAUuBQkCm/JJdU1jagRzKlBXZwI
kn9hZIvnV+hvvqe12FbR/F2uOhlj3a5cS5DcP3OYbh7tlfXJ6IGIO2Icj5Yh7mU83wCSSHOC+yUW
dOoKz6QS09mKGHAZkUZpA/2khzgSKNT860ET1zcRncPyzs6rzlc1umDhupOkit1OkcDMB0LWZ16h
EPzu05umGRqEft9zOcXc7kuGKWwgze0asl8aUFG11kKJDuI8DfcavsWNDCZaFIFoM9R1i+7zWsjK
FYGBFmXc0k0pTGyCpadUZFopS+9dUm4ilSfOhjsnhsAW7+5Fz39cIzPvF8dbJMeSTJqMOOk41E7B
pzMU4TBEmTGPTWcyuRHOjgWdZgOVzZmsukEBixRkH+3jbkUHiOhlOeOylRy2n7l9g4q4aT8eSyVk
A8MOA/6752tw0v6TXulr4CLG/Y9dVikd2/VJ4FIK/+n6SiItBVoze2hsh/CQeHW9fqVOtzwFrepZ
T/IcvjbDJfKGWVGi3c87o1QSCrv1sWrSp75/yoYWV3BRaq4Nr9ZGn+TCwH5OGFGqjRncwDtrJR5S
QMg06mVy1phPD9sWkuvbY7edGpbM6xZxAQmVzKeNJnKIuiABdYgCVtc8uCUrckEWbfLxTr2cKTT1
UEbLrCchYHAhg34G9ha7Y8GJW03Sj0Z9ES7NVLGBrSS/B/w1qoHZYPD6gGO+42X3Ae8Sqokn2zZN
+jKQsrdkHNf7s886+3uUjMH0KU9UQt0DFMHjLzWUl6s5B0wf4Vn0X+4WcuZp7M5o98mP1o2x02VY
dCxwg1RlCigsjXLx1yS2sM2FwpTfbf70QCiodPif2gvqOhP1IS3Bq9X++LqVNGdVyBcjj8J7K3k7
/yzoFfXm5ewuCxqUdDcjI90/mGaymQjdODtwhwsDI8rSu9oRcIsVYPGufK2mtLgZ8Bx+ow9CFWfa
LT5wRTnbX/r7vbghUNi5Vl3HKdKKEwcfEhI8ofw9x8EF0XruQToh/1MQbwc8xo5CjGqHB/QyVV6J
KuFaAsUX3v6YgBKFiE2T+HZlgKD8RcAmhfw6BT1LFJsYJmZ/faPT2iSW1aIK8Qp/b8n3jFMXits8
3NaxTDDwV7iqKJ6Haa7vyoP6Q1IhjEzh1jQAAmZz9E2CO3usTOvCod31avKFMN24sZam8EYX38aN
wCi8JnJTFdMcKN+AraOKd3wJclCKjVeqrb3p23cg83c79dvc73cO88RwosggmCfvpzj01i0tzxhS
EWfmuV4/J00+RZoSpChJtG5LLlstUqE8ppffTd9Q4wQphjrf+KbJcgDqf1Ozs3oy9fIUpl/a0XfM
Zv1n9J34F5mYfahDicN6b+sHGVQH6OjyGq/C5BDDHhurWqn2BRsCjbVFRFT3SliY/5hH+NzV3fph
EUrBoT+48RTBn8Mebje7oiVxu/jpi2aI3BgkNmf+HrFs0/xcwEQ9Mo+WTHRG6VQ7hWOvh+6s5ru/
ISgXKcx+3n8m3JKHgLDcLx/ekS6nZZM8HLLlkG5SjkR5aE1O8ICA+o6Z/tvi78xvw/zsSu857k3d
WfK06b/bPrflzNWKo63ZJFvMbWGfSzYfvC7VHWDibjjT604tlE5VaH8S5/yLqHOyGfJdPwaoR405
wUM3lik63WBCsgP4w/4hieaJxCeJDSY4olqsuPqKGKc3uwmVOUtdx11D5y1F1Zn+YfytAkZxtMJP
BYNBjdl6SSS9jBlhEa4EvvybHIyiuAyy4WNOE4OQUIz0zgMaWVHV1Le/KiMczbZXX7UhyGxaMmlj
z0BdVNTSw25x5z4dnhPHO7sP4hy/jWs9Qui+lVeKcY+hZAoe+ZaqPZDStlZdRZobSHE6L92ex9nt
5s0sIvUF8BrlA+H25ZM9e11yg26yYrOrEpembDbQSjEgZq2M4NUBbB5PaXkYALyLFEA0YsFSWYSX
MaR9Bnluq/xpboDHdVrQwH8aYvFqjEJe3XLddHPelrv4KsgpEpXbKQNW1v5ExZUNSB8pSXeDFo5m
PUBiTQ7l3I6MBGEpqHVJ11aLZoDg/kPKbsevrlbfjwVo29bb07i2xNw5lpv6v52bm+YBl8I6P9ki
6SBcP5pB/FShEKN6vMMAhLKwVqYh+ZhkZ43k5X6Npy/cN+w5HM3/RPhIuIAOBMDpC6xotZYvvQqi
rNRSItKJVol0qqqJgnNRaqZCen1LkA3gPjl10HI12G3tKoAQuaPSIpN4OUC/FRxKL+2UrxWoOt0e
bL3KRyPZAs85rkpE5XO5NJPLupJsdeb027NkiHHp9V9Kh0I5Z3QxNHa9gW+Vxg9gwDSioPqiYCW5
XxZQDXuYpsXICLLFSZizlytktIEdyEKhMKRcxEtWwRrmt2AFExUM5G5VPuGFk4nPWmQv4lk3Tnb3
ZQamDd0zyEG6IGDB3nmqQFRGDgV92ILNQZBMYUW0tsQjt0Nh4oi+mpp37ezVhrMtf+BX0jOdsGTm
n47YxHENXLzuIcR6No6/Q+JZLo3rhZtFui9QwK2oeLzCYkMrQ6a0+xGSFomBvhej4s5vCIt3dr4m
GMDB5qdPuoTynkMY4ilJNp55R69pIPSUmIKtBH4Rd4EH1CRNxaeDITP92wsWd7xAZuwyBXMUehs5
FRnWoPV+RNa9jCfUSZyWb1Kb+TW5T53BxtlNTcdMFG8pEq/+unF5bxCsYgy+OSbz7MJP0pXu9vQB
FVCE8X3oSMGTl5rUoFkFAf7ybDyg8/nb6+/mcVJb1/ftOpVAGxswUTA9d2fkzCZqKMuyWww+jlQQ
yvu9ahIgagl/SRTuxjBwVmZ/zUu1EQZndCJ45EgMO5e6DF4a2DPdTyjab9Zde3kM/UdoDmXJ9STp
s3MsBICXQtEunMl5G9XryIOrBk4SA491tBa/g80FlYhE97YJIzbZYWXPlvpCQ6FsAwmXEIs3QkD7
XUlPjWB3HYKLMhuroYs6JJhi6QSFDFy8KM5upMIXEYtWaiZHaBZQEGRoH67tybRTbzn6JLefo1ya
uUCfPckKvdh3FUJW+Au5Vhi8QcRWT3KftilsuS24vdng5YKlL8l/sGECwXYWG79D/v09lsuJ+LQs
4G030fEiLna1mSzHkCibrB+04t0KqpRTBGmaDNvQzYZfoTkmYMWhKPv+1+R6g+Ln3i9PvRd/etZ2
yIj8fAIhevJS4LUoZsaTzPHtTdQ3xdSeszJRA962e/rfO76pqI0YckS6fazAw+wt6wwbcrMwq8yD
Sdj1iOqlm+qv5w6Lr0sKWFkupsUWsERqqy8zLLfjWDfbRC1zozVSUoEYBBXGrlCNrUsWBi38kz0e
zwHtHLBCjQgL5yfK46nHgvKBztjlvl30VYWlG4HzMK+Ihk/41s8B8xztX+fUlRCPqdoDgobUSn0D
d8sBMENB76SwMAUkArgJPh1LfN02lvoOY52Q/iaA6zKQLe5HgvZkfRFHWiTsCg46oHIqcxUXRlzT
SEv/85NcIa+sVy9s6FTfchLq2NDaDAZZRAfvkvuOSza8Rv81k5FSjanYavtp2/hOEY6jEF2lLr6O
r3Dw55A/7WMK6rRPOiiJWk3K0diXbiHlKNvuzUI0E9P+aiAGGft9tTBhDd1ZuxuhjHp4+ZIULISW
0W2xMkJvFjEzQgarP2Qaxfc6u4fowSfjaeTTzV9gELoavDjGDBmXldPQ/uK7QvZZ3n650JScnfqN
O0gmjLNFX2IxMyqDospuopWCc96m+eVro/0yDxoYg1pFMksmIZA0A9KtD8PO8Xi523Ue56iCLVsN
gLLNpJWbZX1OfhX12kC+ypSWE6jOBfPrhezYKJLrXIySrfhQlz+yncgbTnM1pc1L78FcsR6wDCNl
A8ztqSvLjUC7u/vcDTKbfgTG+CLhx6u/50+hTw89EeddNx0W+ku80tigD38ha1f5At8Yj6/ZxDEd
x6xEj21VxnvZX8REwZercM0Atc1/mOJ/zF7gjRv9PIiCUJoQ0fJR554O4UcE/G2JXsI+Jg3RKU5J
Ura95UC1zxCBGDGj+LBD5fBCa90Ou4mg09hdZaYjL6hJb28GWM9G01YwBPNMRawaUF+WaP3a2rG3
Y8g3UWRxN68jOqLjuNpe2SQBD83O455pCzSP7S1EGzo2i/7eFvMJd1bj9y0k/Z1v7UY6PZ/W8Qtj
58INcM2/jIrpuzIGAVz6wrn2E2s+Oz3hepjfY6549re1L10aL+NOWIgMlczoV/ZzISiDU5ayUNJa
SPZI2LSSx7bgS8pBCS2WgijZzQgwal2hfrXSUHyRPVbI61sErFXl2WPYSK3yWMdqn8cRJh/it0Uu
+l0ngyclvGYmezRdn6brrTDXmuoGuKcXauVDra2vJRHC2GnoVwtTdttEa3xFV75x/QG58wzg+s2N
z68Zi5Ot1HjLhoqshNIqZi1x9ivW99PKcBbzkg+KRAeOGx8DY8NY87YPVVxwh/Ngei0KiO12TFP4
p8uXSX1K4GJBabGPpeo41kqZzneIJTlYqSz9bDsNLl77LnSD6yV8WuiX0x3R/xh0H3IAIxUF3DIM
ft1qQ2cyIAqJGgxS7EbVLwGFFyiqKbM7cEA5c2ni0L06ejr8a8rCkw4gQ1+vjXdeuwnAuSbdjq5K
LXtbLukznR2Mt3Vv+f8o4PRoXv78fgDg3q7jrdx5eETM/Lzys8N6hZRfOL+bQr/yWELQwQOuD2Re
JovMZq8N73duWzDqenUZzpFM1vplA9fxkcqDwsFKqPoJWtLetc8xDQf/lP2zFU+WI+UIPYcyaxg0
SFqVLTqgxRsnfUGkbFSEZiMkvoXw9+PldEdHYhM+gKk0AFYgdGCHc7VEUK4f1fK0u5umayHeSFVK
Z2nF4EjWhg7ftUIsypijgO053DxHXsuYKFc9Nyac34mPkvP7YhcxjzCFyyUqvrORps8BA5yRGGpR
yFAgxCC6kyw8RscPOTjo7XVUQCaI5NCUfSgaJQQ/XP1EMNoPma+xSTWEvF5vFomBz+dzfo9dvu2o
gf1ouwDFXylH+s4geQlFvrlxPwCRiz3UG/S2k2YJVgn5kaLxsA7w/CubX62zeERHSz0YDv7B90+J
6nxVqXhfSrN01Y/SaPQFD15P3e5fAwZmYQGEyIlvYWNzz1jVrDMkKcq24Ndxq+sQtbBjTRJoJkHO
KlzQJDt8cyXmqtSiXlffpANBgiVq7PZyH6zvOSnl7UhP+nFdrmHFup7HJnHOGTpnlKXP2t9qM5qw
aKKu1FKxTibjqaqRM3D+76LjJ/QiAewh63O/48u13uB4MK7imdmcTdX7FdPAVpTVx7JxIpLsTuun
TRvSMfJi9oqr3hA6CQEHgvfGQsHHO0umkBcbgXEJeHjOjrncUyMNE3N+9irjHc6S5Sb472W1sCXH
BmjSnnLUz3Uq/QE5i58GlVwrUeS531zYXV7dav9pkCI7NVM3v6TKXnJ9Z/zl+Zy6di0xXe9Whhtk
OcGTzRSFrIRrq271jx1P4qnsxcwpuEenASwKapTNfJXtxY0iUC4JZrXIkBiYohAEi9JW3rM5qHS/
EjqucCXbPoYhlBwrulyUWPtRm/eEDvOpf0wTFuYoGIRNSU4P2zQkBz5ZjJ3ry4Y6pxUyh6ly9C+x
O01Qj1waMxiCoNR3gCpiUXkygjM+ArihD7OBTO6x+qmJSlJ3yBTk5ghw7yANCre54fAz2d4wC6fY
OSw4a8EgTdUpkvUjCOp5Ylp5MkZpmjFIA51NrTZkyBazwaDSyIIoyf4jZ+XR6BPLz74kU1fV5Vj6
N3whb+rOkVPgjCol85vXozYJ7HTOs1Vt0JSJYPkDBTuEhNeJmFRrP07KAoyWTvY2K2KZlWuzhGbL
ZAZbH7/LeowNxZZlIw7O32MWd8KBtu5f2k/8PEz8vxZp3IaUR4yV+aWWjdX2VLeAQaGj5T2yfKFj
i3wBOS//d3uIKaNl4W+BPezq1WlZJQOoy9STlKBzlb1LR7uDbsPlsO0JGtEBOB/5X0webd7mGW6Q
IC19IWQ609HqL03yPD9DdydXXFoyCYLWnlO3HCmpKzGdSt8pGVsotilF/nEZ32v5pG0OmgXKQItS
mlQQKUnP/VDhkLksQeYMu/cKwwrO9TSfJHzehZKxLvyRQPa7HrlNa5gyRc/toJnVRyTvr4hB0LAk
asc8mq0h6bXr+ldkg72G/j4uF/qEVZIdxfI9IOp4omEhbLR4/KZxXmj/qXyUpaB/6HNiGEbUknc4
Gd/JelGBXpeDX5j34IbHjfkM6P2RfuwVNKbCb8t+RPGPx7rzPyAmPHXFEcUWUgmzNHm/8eVPhNdO
BMbaMl/TcdQC1Rx0TRomaFaaP/o/BVzRo1fHNw+uAlcPDnHFQ4NC8BPGd2mIzyO2+I31usZOkMfu
+SYyP5i7hMFg2K9pl8/kUvus6/Dor7eNnopDRW+Dpxh9A4TSVKuh33aObT0g/4gZpkQB4XMk/gsO
fRJD0gz3+SiJNIVRaML170iKWPi+U3VJg63i72mo4PUVMpNP5FVoq0BxKFd6doaQ94TafMihivRN
gJaQ01sRuxVgC5X+Z5VRlAFSea0JIVNXd2ORaT6UZFrsLKdAAYvlVx2Zy7m7klkOEFhsVfvsSP2S
UawbMab7QjSqdQbLYx5+ck++pNT9i4uFuK3gKt520kVzb2o7X8gBIG/pRbXvdOFoyHhyvhxONnRi
EjSScflEbhrM90Ny/ILArp7qgERZ32USKrkxlfr7lM9oqJzmLyAJEN80f9Rx4ID0d5zRknVgbjsA
7Rg/icl4WVRAg6m/z+IplevbTJg/hNH0E5KR5YoNTchJt+VPw2nVYFf+zsbtSMI7wZ+iLDQoYC3k
SoBBIx0HrW6A4cEf+H68FsxJ/SrkNGm+owRfxtZbiLHPGwy4gTj/JxTSlcgob/6xA9rtbCYIcHQB
A4dlqn9A3A/dWWmrWDtJ0P7D03RmzJcp1MzKOhBbmBlTB0SlPLVza4BdFXFMAgTvQueuzizvmySw
0uaDsp0w46dpztdLG9yhoxMl7s75Nqedw8EFU7H/nEQiVFD4cxb/nUzHkhZpgyXcVeebrg1Idc6Q
1mmuK/ayxRfTl9TiyFpwzTBESeaK57jMATkj2wTXKDJzKbmogQgPVCMXWCeBqnxcBQ7Yx2mnDL5d
bEc9MCfJqVm8P6l1CBtBx/wCjT8PDsh5N+QxLq3JNxqy/5QXHcmuUA4EnR7fq2ePqxZQ13vy+xvx
RrWRtnnwEu94UHNhPjqJJeDhN57koKA6ptA5hP0ZP31/3irPt2GC0UJhDPkj7fYxTDCKAPsjCPhg
C9lJugyGr7vxTjvOkhz9Qtxy5EY/D04y+pcOIzcRyLhzSaxZC7S7IGB7dC0TtOXOC8o8J2dALdBe
yoo/TPf/ikKStARaOM0m7ERXPbYKjcuA0GDzC9MIh5TKR8KIgjQ56lfa+2qofFqTHA5Vhgfr4LEm
+qEZ4on4jVBmzUDAbiB8Ac0HIcVjEAJ9ZtVDkcur1cQLejErpfukToVpUNZZ7CowkrQT9wYJh4IX
FjrO1jZBfL+7C883JJ6cdSk+bv/cwj+ttZa3Ckg4lXH4BB+Gga1SLAjsDbD5YE5BAg6P+af2t2P0
Z7Rod8LAMmVNEuvfBd6J/upux/IEPXPoVWp4q/mHUL/uqIHch0s3cHeXm1UHP/f1XeM3WM5dgBK5
+C1u6JsWs3D9RL/ZCHmk2Pz7uLYM7yy2vw4TDwV0emFAtd9aKWsLZWocZh/QqSt/z4HYcaVKolEc
TC9s8QtvPFtG6PD0UqvA04VEAMka8Ca+GsBkHf49KsqDz3zficR6uyUopE+Oxx4QXQZ41Vbn+kDu
WjSVkTRZVkAXt7EZbML4BbZKVwXP8A5tGgPeAFxICIwH6b0dVyPZ4y4hewmqc3Lh9SJiV7l2NeQg
BhccFZNh2xCkyfF2vZHFUL6S5h9Wb35IcRuXNDmC705UkY0hXvFXfShtwtCz/S8TeiZcpCPSFlMi
shHFL0hiZpUdMhIFX9/HhQU2WaNRv+2JWonUzDHh92g/8uv4rvfG3zDQKJ17SpvsVVrdOqEX7OSY
Io4f/WEXPP/GBeY+0b90UjXiG/ZFmxXLi7UAGGME9Blby71eYMTgQAauI9jT5y22jxkwdwxCxIjN
D6bfv6Uiwq/HPv3VhHSVqJDpUVjUIBEiK97EfwCA+n9L+coAaaCPpSubayO10n5+OMkynSpp8koH
1D23UZkVSFZ5dT35V8WYdO4cVEHYdDYRkPBvgeQUUvySJgRMiZcOOOO/mFLXHKVzQX9zaKpqeDv4
19nKYgcu+0DwPHt7FGETZoLjgwwmW/TQztt+oiPSi+htl4rIOTEjSOej/xzGNTpOIBti6l1ZNuYU
L/Im8O5rmBeJk9ywzWJ4LhrQM65F5S+n2bxpBtXv+t4sYxXuL26J1QlgN2rLcl9Almxgy7yNjPih
LGsvM/YojvPczkhSDfCEs4y8M0W7cCCc2hrLZzSe2JoZqYi1vzjXiIrmlC2fNfXc1HJ7QWkUvIZu
cgVnYHOJMxd/BNcZIBj2pcNgjhgKecuT6RaqNhQiRYzWAf3atn5LPyxFsyhUUuF55h/K2n9l2SI/
hlWJu0xBgSoOhXhIfy7jsG8Pz85iQ/GFJrS+X0DGbF5SHOUVuca6H9kpthbOdo323yOkyOUmMbpR
3BLCr6gM2rbKwJgX4LOblt+z6fR/ylwg65oGSCBVEv4XZ09h2BT4sR0Bb7OM3CS0l5ySSGuLAK0K
rCflSCKbt5Ew56AFh7uwUEmf7r/r8Eexk6bkcCwYuXF4oCuZkJw2XVkcVGr3rA1bokC6Pgy8XrHn
g7nJXKjzqvc1g79Aw6xvOmnMi6qbESX1Eap/Eqi1+YmZQzJe5bvmhduEU+s8FEyX1DUSGLkkAn1q
NHWgb6Gpq+gPSbalCCkad8MUWK/d4g3ncP0jVPI9+ZJu2BIhgBT9rBDpH/llEjfLMvQtJnJtIadT
EbgT7k+orOqPqKEa+VWEZYGs8dCyG2E6gMQmHTp/2AS1WNKVflq4cV8qFxKlAMWEd2FqZjLfE9dm
N+028pejQhlV1WieUnM6U1IUnX4ReRmxayNhx4TWVFbRx1m3Jo/sbK40q/vd1hjrHWZooi7U+tAu
mn6XB5o7GnboyhbRwmxFkVHpvFfu83jfI1aJzd8K2n1FS5XEgj/pXgRpGiK2vvAXOJOqkxnGOyKl
1DRycDZRNismTPK4DpbEz+hKk7PCLNpI9wz2jKWhv8VQFjh23K0QFnvwcSSpK9zfjpy6rLGq7sAA
cTazvqGfCEbn0K8rHGQDJU0OCJGYNVavpsJq/OYAFJUim61XmQSmom+ok7EwaiVnC3hrZf5mM9dD
FDi+q2X5b+Sos7fslRPac9QAaVyZwq4hSRNj8Oj/49OjAukDHcyZj+ohT8jww+YhWZ/5chkgvXoH
YBuoBmNErbBQXccHUhxD2VVkb1IAyS7awKgQGC4pYr9dpAmoaTAH7exa5y9lJgVb9wILq2RjFFwI
JKg75/v3PqCKNm93KSGifC98tViP0XW8vuYYbon5V4kGF8LkrDXQ2tTSZ2OXiwGd3RZKm7JESgjj
Vu9/dfP9qlkUQIy/EgK5qRE40R6TceOfk5zhAuJc4/wWHDOPsfhGiPpnH+HxFNuGBYNur2mmz4yk
azkgJMZtKEid7BE3KhKYgQ/kP/yVmszGvUGktZgU0dJmy338OhMyNRhSDcRmUlVuSP8AB/9ZKT1u
UQyrD3CIvBz55TDbOkIxoHzUq/G1kSeY9njCetZbq29f/vASbarBwQ8HgaGlTkyVnmCJZttBCtps
yuq4vXRe7Ih/SVuH/0PFXV3YgBvPW8sPC893aA2z+IVG17xJQJw23IdkyI5wWUl6oGrVP0Vkdn68
2zVIpcBxtk3KTZXK7YoyoTkD4NpvCOiSZlm35QumI1wzpEZ/EpZtQK3UD3Pxg6iUQzTRrM7Hz1DY
E+6BB3oll8Si0UX0ITaiah0p7dF/62lcareIAdaB0V4Z/D+AfyDbOhbMDIWcbsxbzecQRb5NIIQ5
TkTx07+N33YAKYAwDH2JrtVMQaRFi52SFoIdyu+v4Srm/4F5aP3hV+adD4zyDS5Ma2J0zVjPXb5g
sbv7QXObnhG9Xl6xeqjOvxV4sbWw+1+ijZQDv0gMegtvM0/UIvrCVAgsqEw//k75WiRyO2TKYX9+
2eRJvuGpClpw5XsW8MaGpcwsLhUf1vggi7V+qIbHG6gBuL0TMvEp4tfbD5xKiwJub4ADV9LBgf2l
3UyywsFSY76qSqVxjL/dh2Nv/9ljqMdnUdZXvmSOwtj7WhRpGcC/1vJnT7O+Hr4Yphl4Iwlk18Yd
C7vdx8SBR4mh9AcrV3s6oY7WSNJJIlpD3mVyppuotd0qr8umcVF1xM/eIp7Rv2Sd6Nv9umwt0OMz
EKN9tjNu5zC+86i69rEb2mhx0MAgGUKtB8h4SBBpxgxddmzqPVfGlHK8m0ZApIu3tjdaDOd/AntO
xPT3ueHH/7ZTJRbuXM+qXdvhJSDG31RdNzzjUhsRHLLgk1o/xwjhxBtBbYioxbJCHx929UGPCTy8
CKql/AIaoHRToDYJeiNapjagH09baAWt27ubdq/XiBbJOhf60F8i6+pQYZsHACRg8K4O6rmGjAgv
Pjjg5EZHkZJBvsM0FHp7SDz2vRqRHy2ZRQTdUpXuwJez37tcFwszEj6gXEKbqaraC1B4DRCN35x0
T7q6IJXHvwezdech8HrEjmLf2pCD4RF7nmB9t4oR7+RX8S2FnMbf1ZhFevf80Hm0mbI2Rs4ggzBG
n2YxCUWKfjtXjizyuIX5UvcrkHG9TK3TVv4iCCep+0n5GAuhsU4nHkZCGTiQ7ai5Y5p//THNbHeo
Mp5StGyOUqwRVXMgc7/s/TLVQOYS5HApsxuo2w8FNOmTyQO8ls7LNq9+N1deMno3wEtkIc24gzv9
ULma4mgbIZRQj+MI6+JWVSA4uUvqqqKOssplXZDkZMTNeIrU64bNiid+MsiNd8ag2dBNADXrcRzN
Ocw+GsBn312aoCVJJwRayjQBAoN5hIvr7q4RancU1pfbIBeFB8I7lFxcC+Ogx53ZVCGcDkFjfwfK
bPC5fOpaL7bQo5NUrESzqmLHX3+L7m6RYe4JSprvISL/RGK0YvFO8MT24o0BRvz7QS5rqewgcurR
g22BK2TgiWbPwAIJgWiJ9FZWwBtKrr+bZQqqH71GsaYuJOi8akEHs6KxgROWiBPwdNvmoycts2SV
rwhlHfrHdoKnHvlIhz2HJbvoOoK1toTHVq2Zy/qXGZSHvzSHgnQYwnk7fi+O4X9x68FvSMmQcV/J
WM6/xlZia7elbO4Cf+ok4v9BMm4505hDekFwB7BNnCHuGsyGjhCP1E5t4zIfI6kdAsKCwmO4AT5s
GhTc08zcqzTvRPHuvQq8a4exKyyzO5k3D8NDPYf7E013SE67Ap48lDldGgFqZzOJPF5ip4QYYWLf
Cv4A3ZdH7dOjQXxzh2W/iAbDBkhPL9FJKcCMaq2lEECBb5EsOhJUl+uDICQspE3VmQdqG0Msgm8C
anJG+PkXEW5xZXaaXA/4Toq8RRy1p/DQ3Wzok5VbdSu7k6693iOsDGLoTvukibWPpPSCA+N0/Qao
Yb39tSBM3seMXlsdq/BbqyGoWItt3GQPp4PqMcNyeN74Ha5hdrTyDAuOIFR4CRbM/Gw2mDzq6FpL
tS4iJ9BMBcA6Eq555DPX6fbuthW7XwtN4n0nd4rXWuhuWYrGv0SuBhAAb1XRNei18NTyXdn1vcjX
yZL6JQSE/utmEu3jJbU9XfD+ucPja/rPWjamsH3L/egJZEHHnTsV4eju+1htJ9sNd6e1bHeii+iQ
9CoHwY7aKyxPG0ugP+ArrFwg932eyS5NR7Hkb+GKEwVrk1ew/rlbODybVdYS+uAf9Z6sAMLz1e+e
97BpT826U7D5KYoT1SGyPJOyqU5/HmlT5Oqg6GPK+YH5N5dSA8royrBZQ4POuuagBuQEu1PJ33o6
+EKA+BKMYJoErWTi3/QSwJ1bktIoN7gPrFGqYihfI57XM7zZ3NPP/yEinT5kRb3H81nBaVmH59hS
Ycg+anK/uKVbDWdwqulGFSVR0ELOaKZrvnve9LDzzFbo2c8H1E6n5Ki/xPKDCTXjY+HsCQbd6moM
3tzo7BL5T9SDkyTyyqmbatSL6hHBmtc/E4xha5bKkToFisj1Va8Oxax5A3ElCBM9rjnDmi6tsEyX
SAaSrkCd+Sj8r7V2A8DVEqksKyzg3aI4Du9oKJ9Q6Ai/1wYB3jD/hM13Zm3zvrnEhuO5sp1ilc/x
1YWzVMKanK891rJ6Qwgjw0jWGnBxLdq/jTPopdnouFi0PabMyI9HOHkC8UddzqNJonprFj4aoQ8C
T2Ome3eLb1+qLi33uN7+RyEHfueTiE2aqbuE2bswD5+EHTF16bTncHkgoxrRKzPujFHfK0N6D/n/
rCiN0oa0b3GPx+3ZNHpqF3WJr1eFAglOUtYuD6sSWbJoUButNTA/rFw36ZB1SMFCLInpWy/H1jOT
z0+VgO6Em3EvS/R7UnCI6R9Qjy+ZcVE0FrggTcP9nTrq0+W4tinQxyjHhKN7LtQKJ7F/ZvHsn8nl
X3PaHb+/BA2DjTB1hMkU28LgbGkFq61ffMiYVoQhsv7Mf385TKcygrNMTJM4bFRUeBLKNDWFwRQL
Lof0vSLAJzYCnnI2Zjb5ME2WVzKunhNmB+LyU5tXZbPMl7ZPfaoEx2rjFIV3d8Y72PWGuVMzOv5n
XernScoFGVGtASPzd3uXqIwsCe0IWwZEvz/cBC4hwPO/FXVzg78ZNqrEKF8lp83m2RLuewyRzAmV
neTEdJisnq6Xmea8ivr8EDNg1HH7AnD4eiNWcL7nuDJCpfgEdiIR6P1lOXgi28SelspPSviKDLZg
vqGwNsGQXu2tUnzSfmoJPau1A/3Grw4HdhvgoL6mkvl2DSudVDhAEtjxonilefU0u7l/ROTaw+xF
/JgtAu/eZm2GgByLzLyWY1qggswm+EfCSUktg7LgyEP1IE8iUgRR6ZoUm8tGlVIbsVBlM/x/mlIn
+Do062A0YxnsCb2DBvcQv3E2fcsHu6bUYC7T5uOXqtujpu+QnVjihalCnAaBB8zUJ+SjLDh9cq6X
P4osLhut43tRt/dcoaUb9Lr62WdRhGY58sAwe+z1hP9KmX3NGdFgroTy6ao/y+kMjX4u762rn3y4
1J7KPRt1rutOnzJ4hVgA2wIRB/zx9WhNn7TFdRZ7V4m0s0u0Aj4rO2OOnbV5rXxLSvQ1EotS0XmP
KBI+cfYXYtEiZtRPHIvOMjR2yL4aBQJpfwQyX9xlf5a4NOl8UTHokdFPncZoRwlwoiyOumo8dOYm
VfC6rLyQCUQU7+shLElPCRsYSeKZBaNZkjUyOWBoCPaVxCaOOH35EJ3WCk/D99UBUl3jgORRTY2A
c9eTfJlMAEcsp3P4jWUJ3Zog0C6yP22M58siF/3vQ76Wc3M2slwuYqDwax9mH/9dh0eAQfQyI1RX
6g5yaZe+yb7hhk1XM+2exhVDHEugFTaf1b0REeKcnlnn2bxPhDuW3EGGSMlECF9SPmsFiEedzX5+
yHSSwrA4baa/VYCv36etjEGNgDW85yZUZ/cMn9hMJCEaIqK8G9T/A+pIwcr1LgG1XG9DgA55BQi7
TqGZIC4RBHC7dQqOmTu8US4hVvnH2ASWg+Jtl0Fkgtu8kRjEpwV0g0KVvlxr5L9ovG6HhgHSBxD7
omsXyBfjmdMm6aEUBO5j67kL9QLQXnGDGGgj1yskWiJeNyhVYTFkch2xhZLO642gmZDhJHgL+NEx
tBHbR83bOeb3O4jWGbY1xDod5ojn1OgkX0CKRAwNRzqXjlQBPCTNqfexB4yYtUMeAcE0gRiRX0o5
ocDN8FXM6G2ZdK/sI/Z4U/bJ8RTqr2bDqf3BF3b7icDk9Qy93v+ktZX3rMw3Pu1bUH1D6WyK3JCK
e9GsOhCyH5fjGbIRxCseCEW5ID7V2kZKM3uNHIFzP3gsJLCyYzZmTbOYxCemfCDPARGpS1goqGv2
S+uf3/h7+1M2webQAjrCkM5k/DLGoBTcSjAtE7UoHFVaJ6qcRxbTG6facfTBCcxLkHnM3DJ1QHvu
DIgoxPk2ZQpwT0zmk0MhjEWMYYUyHk4cbSi22JfnFxsXhaIknALf7rafE1pk44fFMLcC8zh3yhHI
njvBRAx5HZ9eBMNSnLKSACGyEDMfvcafqt/Xq9px98h7uIohVdNXwXZKDY5EU8ItkisrbsCQOPH7
IZKbvClbzA+jaQ+BUl9C5pDx7eO70FthnW9FHuc+whr+c5Jvv7dq6t77nl2Vavn9F4Lppv+ohUrH
S12sjX6DFra+yiCt0u+dy5tjBKwYVgz0yZo8Y+CvqKzocIOaNNIBLlksORAJPxR7HolGc2kXpoWN
XAr7/DPNgnPwUZP44S5LaPu/cjzv4MC+lgKCHUrwzlfXCHBql9EClb6US9TmklSLYwJ0l1zDNnFQ
tGWFdx/PzqMsca8BxOodeqA6c1XUpRO4/8H+S6kwAeISY9CMyrezN1fty7H7eJ+gab3K/JKSo9qe
h2Eqiou21ECr+6jDNC9A7/6S+p5RYGTedVILw0Y0uvBsrpd4Cg0ngEaKrfdpVPqmxI4MFFjcB9b1
Fr4b3QezEyrmL0lJJ1Y53S1CU5XP34DqnqKjWnGIv16yWY1qCoYXccE92GJV4Rha72UThfH9aTfV
ETx2uBdc6zzJ639xw4u4OIH4pX7YS5HPa2nlSxcoaj4rYCIw9JcHk92sFHWET8QUBlPpV3cVZcNA
mK/NO57Jl52mjseqFkF81Se7RYTI5n7/09e65Ejtu4BGSkEakSFfOIR5OPt44++pVvfMlgDCn5kn
d/ZDns4+tq29C6JzsLPdN67Vm5ctYso7xDCsoXfQgnHtR8AwRim3VTWxOdwCCOfac9CQ0qKftyCR
t4JKPnUZGjHxiTLmeBUkKoRQxMy7zkLL1dh3UhQKnD3X07nOALIF6kbN55WW7Lsq5A/yJbjBLA7j
8tdbnX34hvvkPkrsia+ovLQYCBGQHIClxjgte18b/oeYGbFw5oeEnE7+H3TmSKGpNYp9d9fdPoMt
UDZ4PWeCeY1KvP92/7yEAguNd5J5MKVJAIh2EcdFLIx5uMT+tFs2LUj2bg4tXP3ASENY7vlz5GmD
dJoi3hm4BBjjilygzeCv+qjyNEeHy3FbenIxGtFtuLgWTpxlrvpiImnBzmuSpjmA2DXxAvRxuepE
u5UOPYxTOXPdXPc+QvUG8UdujQOIsfJTLzPKjJrAJLYlzCqLOa7xDeSVKArIy/UB9DZgT5uVGQjQ
XebSDNQ4ojRq/Uo5pxDRJrDnIxD1avEEsucYr/X8EK+WlLCiW9aY+XXHzLm4q5+fTxd4HfZiaDno
NcJ6jskjKF8I4pOLQsrCxUnc9Z2vlpWQ1udOsitNlpTrdZhZp83qWrS6ZHuElLF7zG/YZ8V4ywmd
cconkorFrj2x94S5l+6nU9A2MHxpX4cE17r28hglv/pYgCCA7IxMoiszeD9UOuCdihETZqYDqs22
vt2p4ikWk8FZb8Y+TCKNd1ECvjSUDFPzuDVcHd5l8i8tKb0gWLpvoPa3txYCo1PiZHvlLvEyaArT
RZg8EoHP8mDzPVhXTk6HEEq9biUxKUAYL5ysp36JZbk/TcVO2CqOA16Cbc0KwCa58Sr4xuTxAUEo
maOt9ngS4NaCtQT1WNtES7mBC76rGJPR5rGjn4/hAYIuUXSIPlUroibf6eLuIuBDvJoRcEgLxLQb
wnrTBlphAi7jNu6R65Qa+Hqdrq/eHlNFoFaLYkFsx8ksuiUVfuW2GCBDG269Gv40gZQeIJqf4iv6
hhaJpxrCQOfMTtITPkrvuYJdSCygfRKtT40R434zcaeAgcFq5Ljuv39EVGdwFMQLSDMtcd5VfbpT
RVHHlkqRcQWiPXzzdC2IDhGTigneA+WFRHO41ETKFNFYuLnlGR6OBThsZXuA3LPDvUrsOCjiIg3T
Xfb7XXDPlWyl1mTAhnbi7dILtiKTJtJsx2+c/mNErSa0A7a43mzh0tlv/xs9BwkAbI9HcolznZqm
Eun+qk+LCv0ItqXPkMktXNQu2/8iCQ7XPhGhKr1ERdj1r4ku6vsI9cabSNqTcwiPfRmOQxoyHWK+
3xsLF1R32xO2
`protect end_protected

