module prim_lfsr (
	clk_i,
	rst_ni,
	seed_en_i,
	seed_i,
	lfsr_en_i,
	entropy_i,
	state_o
);
	reg _sv2v_0;
	parameter LfsrType = "GAL_XOR";
	parameter [31:0] LfsrDw = 32;
	localparam [31:0] LfsrIdxDw = $clog2(LfsrDw);
	parameter [31:0] EntropyDw = 8;
	parameter [31:0] StateOutDw = 8;
	function automatic signed [LfsrDw - 1:0] sv2v_cast_C2EBB_signed;
		input reg signed [LfsrDw - 1:0] inp;
		sv2v_cast_C2EBB_signed = inp;
	endfunction
	parameter [LfsrDw - 1:0] DefaultSeed = sv2v_cast_C2EBB_signed(1);
	parameter [LfsrDw - 1:0] CustomCoeffs = 1'sb0;
	parameter [0:0] StatePermEn = 1'b0;
	parameter [(LfsrDw * LfsrIdxDw) - 1:0] StatePerm = 1'sb0;
	parameter [0:0] MaxLenSVA = 1'b1;
	parameter [0:0] LockupSVA = 1'b1;
	parameter [0:0] ExtSeedSVA = 1'b1;
	parameter [0:0] NonLinearOut = 1'b0;
	input clk_i;
	input rst_ni;
	input seed_en_i;
	input [LfsrDw - 1:0] seed_i;
	input lfsr_en_i;
	input [EntropyDw - 1:0] entropy_i;
	output wire [StateOutDw - 1:0] state_o;
	localparam [31:0] LUT_OFF = 3;
	localparam [27887:0] LFSR_COEFFS = 27888'h600000000000000000000000000000000000000000c0000000000000000000000000000000000000000140000000000000000000000000000000000000000300000000000000000000000000000000000000000600000000000000000000000000000000000000000b800000000000000000000000000000000000000011000000000000000000000000000000000000000024000000000000000000000000000000000000000050000000000000000000000000000000000000000082900000000000000000000000000000000000000100d00000000000000000000000000000000000000201500000000000000000000000000000000000000600000000000000000000000000000000000000000d008000000000000000000000000000000000000012000000000000000000000000000000000000000020400000000000000000000000000000000000000040023000000000000000000000000000000000000090000000000000000000000000000000000000000140000000000000000000000000000000000000000300000000000000000000000000000000000000000420000000000000000000000000000000000000000e1000000000000000000000000000000000000000120000000000000000000000000000000000000000200002300000000000000000000000000000000000400001300000000000000000000000000000000000900000000000000000000000000000000000000001400000000000000000000000000000000000000002000002900000000000000000000000000000000004800000000000000000000000000000000000000008020000300000000000000000000000000000000010008000000000000000000000000000000000000020400000300000000000000000000000000000000050000000000000000000000000000000000000000080100000000000000000000000000000000000000100000001f00000000000000000000000000000000200000003100000000000000000000000000000000440000000000000000000000000000000000000000a0001400000000000000000000000000000000000120000000000000000000000000000000000000000300000c00000000000000000000000000000000000630000000000000000000000000000000000000000c00000300000000000000000000000000000000001b0000000000000000000000000000000000000000300003000000000000000000000000000000000000420000000000000000000000000000000000000000c00000180000000000000000000000000000000001008000000000000000000000000000000000000003000000c00000000000000000000000000000000006000c000000000000000000000000000000000000090000000000000000000000000000000000000000180030000000000000000000000000000000000000300000000300000000000000000000000000000000400000400000000000000000000000000000000000c0000600000000000000000000000000000000000102000000000000000000000000000000000000000200004000000000000000000000000000000000000600003000000000000000000000000000000000000c0000000000000000000000000000000000000000180030000000000000000000000000000000000000300000000000003000000000000000000000000000600000000000000000000000000000000000000000d80000000000000000000000000000000000000001000040000000000000000000000000000000000003018000000000000000000000000000000000000006030000000000000000000000000000000000000008040000000000000000000000000000000000000014000002800000000000000000000000000000000030006000000000000000000000000000000000000041000000000000000000000000000000000000000082000000000104000000000000000000000000000100000080000000000000000000000000000000000300060000000000000000000000000000000000000601800000000000000000000000000000000000000c0000000180000000000000000000000000000000180000006000000000000000000000000000000000300006000000000000000000000000000000000000402000000000000000000000000000000000000000c000000006000000000000000000000000000000011000000000000000000000000000000000000000024000000048000000000000000000000000000000060000000000300000000000000000000000000000080040000000000000000000000000000000000000180000030000000000000000000000000000000000300300000000000000000000000000000000000000400200000000000000000000000000000000000000c000000000000000018000000000000000000000010000000004000000000000000000000000000000030000c000000000000000000000000000000000000600000000000000000000c00000000000000000000c00c0000000000000000000000000000000000000140000000000000000000000000000000000000000200001000000000000000000000000000000000000400800000000000000000000000000000000000000a00000000001400000000000000000000000000001040000000000000000000000000000000000000002004000000000000000000000000000000000000005000000000028000000000000000000000000000008000000004000000000000000000000000000000018600000000000000000000000000000000000000030000000000000000c000000000000000000000000402000000000000000000000000000000000000000c03000000000000000000000000000000000000001000100000000000000000000000000000000000002000400000000000000000000000000000000000005000000000000000a000000000000000000000000080000001000000000000000000000000000000000186000000000000000000000000000000000000000300300000000000000000000000000000000000000401000000000000000000000000000000000000000a0000000001400000000000000000000000000000100800000000000000000000000000000000000000300000000000000000001800000000000000000000600180000000000000000000000000000000000000c00000000000000003000000000000000000000001400050000000000000000000000000000000000002000000010000000000000000000000000000000004040000000000000000000000000000000000000008100000000000000000000000001020000000000010000400000000000000000000000000000000000030000000000000060000000000000000000000000050000000000000000000000000000000000000000080000000040000000000000000000000000000000180000000000000000000000000300000000000000300000000300000000000000000000000000000000600000000000000000000000000000000000000000a0000014000000000000000000000000000000000108000000000000000000000000000000000000000240000000000000000000000000000000000000000600000000000c0000000000000000000000000000080000004000000000000000000000000000000000180000000000030000000000000000000000000000200000000000001000000000000000000000000000400800000000000000000000000000000000000000c00000000000000000000000000000060000000001000008000000000000000000000000000000000003060000000000000000000000000000000000000004a400000000000000000000000000000000000000080000004000000000000000000000000000000000180000003000000000000000000000000000000000200001000000000000000000000000000000000000600006000000000000000000000000000000000000c0000000000000000600000000000000000000000100000000000010000000000000000000000000000300000000000000600000000000000000000000000600000000300000000000000000000000000000000800000100000000000000000000000000000000001800000000000000000000000000c0000000000000200000000000010000000000000000000000000000480000000000000000000000000000000000000000c000000000000000600000000000000000000000018000000000000000000000000000000000000000028000000000000000000000000000000500000000060000000c000000000000000000000000000000000c00000000000000000000000000018000000000001800000600000000000000000000000000000000003000000c0000000000000000000000000000000000400000008000000000000000000000000000000000c0003000000000000000000000000000000000000100004000000000000000000000000000000000000300000000000000000000060000000000000000000600000000000000c00000000000000000000000000c00600000000000000000000000000000000000001800000060000000000000000000000000000000003000000000c0000000000000000000000000000000410000000000000000000000000000000000000000a00140000000000000000000000000000000000000;
	wire lockup;
	wire [LfsrDw - 1:0] lfsr_d;
	reg [LfsrDw - 1:0] lfsr_q;
	wire [LfsrDw - 1:0] next_lfsr_state;
	wire [LfsrDw - 1:0] coeffs;
	localparam [LfsrDw - 1:0] DefaultSeedLocal = DefaultSeed;
	function automatic [LfsrDw - 1:0] sv2v_cast_C2EBB;
		input reg [LfsrDw - 1:0] inp;
		sv2v_cast_C2EBB = inp;
	endfunction
	function automatic [63:0] sv2v_cast_64;
		input reg [63:0] inp;
		sv2v_cast_64 = inp;
	endfunction
	generate
		if (sv2v_cast_64(LfsrType) == 64'd20056519619399506) begin : gen_gal_xor
			if (CustomCoeffs > 0) begin : gen_custom
				assign coeffs = CustomCoeffs[LfsrDw - 1:0];
			end
			else begin : gen_lut
				assign coeffs = LFSR_COEFFS[((165 - (LfsrDw - LUT_OFF)) * 168) + (LfsrDw - 1)-:LfsrDw];
			end
			assign next_lfsr_state = (sv2v_cast_C2EBB(entropy_i) ^ ({LfsrDw {lfsr_q[0]}} & coeffs)) ^ (lfsr_q >> 1);
			assign lockup = ~(|lfsr_q);
		end
		else if (sv2v_cast_64(LfsrType) == "FIB_XNOR") begin : gen_fib_xnor
			if (CustomCoeffs > 0) begin : gen_custom
				assign coeffs = CustomCoeffs[LfsrDw - 1:0];
			end
			else begin : gen_lut
				assign coeffs = LFSR_COEFFS[((165 - (LfsrDw - LUT_OFF)) * 168) + (LfsrDw - 1)-:LfsrDw];
			end
			assign next_lfsr_state = sv2v_cast_C2EBB(entropy_i) ^ {lfsr_q[LfsrDw - 2:0], ~(^(lfsr_q & coeffs))};
			assign lockup = &lfsr_q;
		end
		else begin : gen_unknown_type
			assign coeffs = 1'sb0;
			assign next_lfsr_state = 1'sb0;
			assign lockup = 1'b0;
		end
	endgenerate
	assign lfsr_d = (seed_en_i ? seed_i : (lfsr_en_i && lockup ? DefaultSeedLocal : (lfsr_en_i ? next_lfsr_state : lfsr_q)));
	wire [LfsrDw - 1:0] sbox_out;
	localparam [63:0] prim_cipher_pkg_PRINCE_SBOX4 = 64'h4d5e087619ca23fb;
	generate
		if (NonLinearOut) begin : gen_out_non_linear
			localparam signed [31:0] NumSboxes = LfsrDw / 4;
			wire [((4 * NumSboxes) * LfsrIdxDw) - 1:0] matrix_indices;
			genvar _gv_j_1;
			for (_gv_j_1 = 0; _gv_j_1 < LfsrDw; _gv_j_1 = _gv_j_1 + 1) begin : gen_input_idx_map
				localparam j = _gv_j_1;
				assign matrix_indices[(((j / NumSboxes) * NumSboxes) + (j % NumSboxes)) * LfsrIdxDw+:LfsrIdxDw] = j;
			end
			reg [((4 * NumSboxes) * LfsrIdxDw) - 1:0] matrix_rotrev_indices;
			function automatic [(NumSboxes * LfsrIdxDw) - 1:0] lrotcol;
				input reg [(NumSboxes * LfsrIdxDw) - 1:0] col;
				input integer shift;
				reg [(NumSboxes * LfsrIdxDw) - 1:0] out;
				begin
					begin : sv2v_autoblock_1
						reg signed [31:0] k;
						for (k = 0; k < NumSboxes; k = k + 1)
							out[((k + shift) % NumSboxes) * LfsrIdxDw+:LfsrIdxDw] = col[k * LfsrIdxDw+:LfsrIdxDw];
					end
					lrotcol = out;
				end
			endfunction
			function automatic [(NumSboxes * LfsrIdxDw) - 1:0] revcol;
				input reg [(NumSboxes * LfsrIdxDw) - 1:0] col;
				reg [(0 + (NumSboxes * LfsrIdxDw)) - 1:0] _sv2v_strm_45112_inp;
				reg [(0 + (NumSboxes * LfsrIdxDw)) - 1:0] _sv2v_strm_45112_out;
				integer _sv2v_strm_45112_idx;
				begin
					_sv2v_strm_45112_inp = {col};
					for (_sv2v_strm_45112_idx = 0; _sv2v_strm_45112_idx <= ((0 + (NumSboxes * LfsrIdxDw)) - LfsrIdxDw); _sv2v_strm_45112_idx = _sv2v_strm_45112_idx + LfsrIdxDw)
						_sv2v_strm_45112_out[((0 + (NumSboxes * LfsrIdxDw)) - 1) - _sv2v_strm_45112_idx-:LfsrIdxDw] = _sv2v_strm_45112_inp[_sv2v_strm_45112_idx+:LfsrIdxDw];
					if (((0 + (NumSboxes * LfsrIdxDw)) % LfsrIdxDw) > 0)
						_sv2v_strm_45112_out[0+:(0 + (NumSboxes * LfsrIdxDw)) % LfsrIdxDw] = _sv2v_strm_45112_inp[_sv2v_strm_45112_idx+:(0 + (NumSboxes * LfsrIdxDw)) % LfsrIdxDw];
					revcol = ((0 + (NumSboxes * LfsrIdxDw)) <= (NumSboxes * LfsrIdxDw) ? _sv2v_strm_45112_out << ((NumSboxes * LfsrIdxDw) - (0 + (NumSboxes * LfsrIdxDw))) : _sv2v_strm_45112_out >> ((0 + (NumSboxes * LfsrIdxDw)) - (NumSboxes * LfsrIdxDw)));
				end
			endfunction
			always @(*) begin : p_rotrev
				if (_sv2v_0)
					;
				matrix_rotrev_indices[0+:LfsrIdxDw * NumSboxes] = matrix_indices[0+:LfsrIdxDw * NumSboxes];
				matrix_rotrev_indices[LfsrIdxDw * NumSboxes+:LfsrIdxDw * NumSboxes] = lrotcol(matrix_indices[LfsrIdxDw * NumSboxes+:LfsrIdxDw * NumSboxes], NumSboxes / 2);
				matrix_rotrev_indices[LfsrIdxDw * (2 * NumSboxes)+:LfsrIdxDw * NumSboxes] = revcol(matrix_indices[LfsrIdxDw * (2 * NumSboxes)+:LfsrIdxDw * NumSboxes]);
				matrix_rotrev_indices[LfsrIdxDw * (3 * NumSboxes)+:LfsrIdxDw * NumSboxes] = revcol(lrotcol(matrix_indices[LfsrIdxDw * (3 * NumSboxes)+:LfsrIdxDw * NumSboxes], 1));
			end
			wire [(LfsrDw * LfsrIdxDw) - 1:0] sbox_in_indices;
			genvar _gv_k_6;
			for (_gv_k_6 = 0; _gv_k_6 < LfsrDw; _gv_k_6 = _gv_k_6 + 1) begin : gen_reverse_upper
				localparam k = _gv_k_6;
				assign sbox_in_indices[k * LfsrIdxDw+:LfsrIdxDw] = matrix_rotrev_indices[(((k % 4) * NumSboxes) + (k / 4)) * LfsrIdxDw+:LfsrIdxDw];
			end
			genvar _gv_k_7;
			for (_gv_k_7 = 0; _gv_k_7 < NumSboxes; _gv_k_7 = _gv_k_7 + 1) begin : gen_sboxes
				localparam k = _gv_k_7;
				wire [3:0] sbox_in;
				assign sbox_in = {lfsr_q[sbox_in_indices[((k * 4) + 3) * LfsrIdxDw+:LfsrIdxDw]], lfsr_q[sbox_in_indices[((k * 4) + 2) * LfsrIdxDw+:LfsrIdxDw]], lfsr_q[sbox_in_indices[((k * 4) + 1) * LfsrIdxDw+:LfsrIdxDw]], lfsr_q[sbox_in_indices[((k * 4) + 0) * LfsrIdxDw+:LfsrIdxDw]]};
				assign sbox_out[k * 4+:4] = prim_cipher_pkg_PRINCE_SBOX4[sbox_in * 4+:4];
			end
		end
		else begin : gen_out_passthru
			assign sbox_out = lfsr_q;
		end
	endgenerate
	function automatic [StateOutDw - 1:0] sv2v_cast_7F415;
		input reg [StateOutDw - 1:0] inp;
		sv2v_cast_7F415 = inp;
	endfunction
	generate
		if (StatePermEn) begin : gen_state_perm
			genvar _gv_k_8;
			for (_gv_k_8 = 0; _gv_k_8 < StateOutDw; _gv_k_8 = _gv_k_8 + 1) begin : gen_perm_loop
				localparam k = _gv_k_8;
				assign state_o[k] = sbox_out[StatePerm[k * LfsrIdxDw+:LfsrIdxDw]];
			end
			if (LfsrDw > StateOutDw) begin : gen_tieoff_unused
				wire unused_sbox_out;
				assign unused_sbox_out = ^sbox_out;
			end
		end
		else begin : gen_no_state_perm
			assign state_o = sv2v_cast_7F415(sbox_out);
		end
	endgenerate
	always @(posedge clk_i or negedge rst_ni) begin : p_reg
		if (!rst_ni)
			lfsr_q <= DefaultSeedLocal;
		else
			lfsr_q <= lfsr_d;
	end
	initial _sv2v_0 = 0;
endmodule
