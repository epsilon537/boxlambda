`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ekqTGLVeLCGZCJiiSNF+tMyH6RwvcLd0xadQIoYc+Ag7wn9cTT/S0FzABqtmRFpQIv9pKH/qSef+
6oY3VUZJqZ0nVY7tIwaT7CH/eiFvMnGvV7fL34BqrQmLoDvmNEFaor/cgwNiFstMNFoJyXXmp1p+
Ghs7luB53ie2a5UboJPmjRMKe1Sc/YGC1ROCCkIufwwPMlUKlzZRus3K918PFVER+X2rPeTgaR4+
J+tJsdYcqLuw3MFMW/57u6B7RvdP64QHEdMjbXOGubWQOVXCNJdKsUEuO74HSVtZ+ArLRhFNtzDu
MvAvVCdjJNBdFOTPhhfUqYaM0h+zE8W3lOZKcA==
`protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`protect key_block
jSkEK8xaCt+lTeaEsln0Vp6C5yLnd50aZ2jgpuNe6uoF+S/dZHpcfkQj+Dz2T5pG6RdKM/+gUjcs
epcklxJ1xa6gq7b9qUedRmWIcvUzOXrq39F2W7XssoJReYTN4oIin/cb5Qdovn/uwWYM3SPG40Vv
534C4bz1LWASSNx2RpsWqytqMtgrDZq8uEVoQA89ixjL8W6DzYjzXh1ZeFEbj8vPXSUzU4ZROXXU
1Mhlbu09FBAOwJWyN3U/rCcHlqdi3mxME2LL7AkkS6YlMipRNfx/u3BY0V82rTW2Ex/a4mCBBQvT
NBzPtanwdt8YkpQ76xyDzGfbwwKarOEpUwxEkQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
q0EdmEvHyPKr+d698qLC4id46xzK9evjroqwPmVY/YVZh8tF+0uaevOp2Y2+XD18iq2gZMLyk0Ms
pLr8t/sXuQ==
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZE/YQMkoOP/F8+QPEPjohNVTH+DwVdrz8uEHvycuem5Qs0cYOQvmin4eQRWq2QBTqoCXasLoiIga
QjbrSd7Nv+1LMT2j3QMzuem7DhzUwqEv2Nztt/dzw5QjlAoqAcjWXlvxe58tdz82fuXFSV54vShs
duN+nmUPlrpMAG8zSPyup27B2orVQGeAn+QGZM12B3Hvpqr3eWblJIOo1tURo1Z3IR00r8xKuNp6
fhtWa6e2zfNKmx3WO2XkJGWFimgNJlLfscKrfBpzVvFjlCh4hz2ktjafAk6OmD21WgZqS/25AskM
Ya4peXcPKWy+zozb7nVKYwiFekza6uVD//rvKg==
`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k5oRTY6yPss7Z6PyCZwRklbNez4rFduKqSswPxWfnSHiXKJXAnuy6e7QX6kR3AoUgJHFxyn4hEYk
a+Gum7Q4eTASWzXbPHDH1gzOQi9Jo0ipWhqzRA8JTEWWFO3IOLAOLjWsuoeGam2ftFqIlyafyIOt
eRldWnMJbZbdVrMw/Y2OyXMeFR/1/sirqo8FL4zXWdSLtGZN/0ZwMoqNPCJh4GtPMToQS7jXihrh
rc/OG/17rdNMmpwcWc0eaKSKztZTE/Sg2fmDd67dnaxVeduv1q9PyvAwt3lHSs1YWlGHOzcLc+0Z
uChwwj4eWZzUnyE2LWa93FYyd+xzOmTGKXc0Tg==
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JoW7JdY+gPZERN/qVjK1bt5mYxqSnILneY6/ZsLUz3vIUIyJpCfQHDIHMW0tw4AXJbIIdvmedxHJ
iva7MFtw5WbOpbM54rcYZ9tkEC6mHK65Za4N/BVavrNsvYlFa3igWuYnF1p4PVx2C6jugZYyk/rJ
zd89pn2tuH78jCBOXR0=
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q1REQ1VZuBhFwy1v5fnnOV6YUS3qlDoQdFad0k3P/Iq/fxQ7S5ugOyE8Q3C+5TMOUfdHrUCi5C3c
jFtnRGRYlm97X/+3KRp49yCmOYUiyxA0fi97Y2OAMiwQ7bB6LgYkKH28BTe1mDped2Zq1E7agZSC
B7SAa+B99J6yqsVlFjqRy4oldaUnRqD7bheMTczLZmqLSPW2hhutbzqbw8zQ2MYMFo0xfYCZ5fTc
aV2+bxaWBZJzP4EexcqV14tsXQnbIBm0S9GMI9zliP/9bmp38OUUOi4fb/oo0yBco7EVboRk8bdW
WudRaFdm3eYSokQ8B+PKDGcqyMgIbEHjoIluxw==
`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JJHW5baXz+5OLs35TBwcxJBTQWRYAyr064oNN6X/LSDaZAZ1/KPX7eIZ+MwGJ8+4AGDViLaczYLN
wbCZnjoK0TO5lAE6jWTebIsKg8It2+XuE+ISWtolQ272yMWjsG1L/IUIyvhBkrFM7RrnMbFhTEYu
x8RYyjkFAkhBlIqs800Bx0OZLf8aZXyamT2gjiznGruGyZdnvAd2F0q9GH1VfgSuIVvPnBoiKdHq
oNFiKTuIP+uyX90QWdv2AZ6FAy/nGWVcjpVbGtVoAWOvHhiTUqBSz29oTzWDIp5EntXsRjf6zsPi
J3poGNjc1JNQADf8i8mBe7Tr54A0B0awFv9X1g==
`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bIiqDkmm6DX/J/hle4I+HBRjha5QGkkMqCa9zyDt9h3U2VCO4OnSh9FD3neJnjJR02pSwMH0Lxfi
saMSMRjlE8+2GZCR5GScqMMdSjuHPyDQlhZ8ZQi0vug8jlFZMsh3oRJU1ZAK1Uvu1ThtYcdiAj8f
IdbdiKj8Q8ZdtHR1sVg=
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rrUA3IWCjN7ulbmOC0knw0xVonpwOG7AWa2Fwea2ohQN+8rngh2QVoyzbfy289YPfuV0uesPJw/R
g6ejJqpVrr7GgWAmayTPzL4g2661k0vz6D3zf3tyCqpkVDe0CzZkVe1z64jDYRtDIR8sAnj9B53w
PhbhlPOhCc3qXxst+ZJYGq9gbucQZ6etBxwi7FQiLboimAhPrW5whCVdfHKIrsAcGCEt2tVXs2kU
Jk0wO72vy6T/st+EqtTyekLn7qaCP/YbCsdS27Q+B8K9rm8GPNOKUKIYxTURvx9TMP27+zuKzseG
iDCi+3xjYmXpce4V6mjjbDhnwDL1ZojrIuWuEw==
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 206048)
`protect data_block
beUbNnLh9kxjMl7/R1IAtrWd2yTnyWwR1WfaIw4xns/xBAXW70iXb/tMEBvq6vfNNpsN6YpPSZe3
zmN/Nx3h2drPYbwyV5JoL5PnLe4cmePvR8Xwbl4mLR5Uy4hJSC7HT3jOZZlKhOiOi5ubFcESHMqH
d0x30XOobQU5Aad+XWhPRgZz49wqDLEAMyJyQ4kFjXhc2Gjq4I2H45T+4lFZm9D2M4dw/U3ypM9A
r5Dujv1nfl8+x0Z8ulXAnuMdQNFXhotF9Yc+BwgGokef2ct4u//mymPvDkTfEBLygIgFmXzFkmKq
7u6taJGJ8ncqWmIG7aGIiKB04FrWDz2vaGswm9xLVnLRuibuoV0VGAdGwgPOA1ZeosSCdFWMfUgF
fEHc85XnTlRFJElkVzRDC+66+xTAxzT07Gmj3DVaxn7IThogoYJC+s2j+lSJC9bHzbtmP5MxeCF0
UIRfN8b35yA+ZvpE6X222g1wr7U/Sdj9OlOxKByE+078NtnOqERCxS0VgDeN+T1TpZLG54m7+Xf9
yjA2xVao90Wd4qzVBwqbluibmrNRb2OdikVG6nkpLwfhk+woG4P0nTw0SETCez8bZOXtVDhrRwQK
DHYmVaFvYpo7CDPdJ4p8KGQPvGWHu53Nup3wfGZAOVB2gTyZEJFA5aV6PkGRlRELuI5BKL8VzQ1t
TbLNR1YF4/n8dv214prq0Q3NSV06rq+O+fAnX2e7YxcOFvU7dl6ApzHURtCatFt3VjTxzTpfqGzg
xpoGmbLJKkRLWgi7oh9bklRuhFpSktblTcRpaUces24hcYRCaxw/UL2EWu6X7zsLeXn18uNrWE1t
WJjhBKfco2kcSzPI2xmXGbiFaud58p2tiV84zJNlkhlXr2qYs5ojVBpLOsxpzYv8KtZbFQ60sRc6
WL+70JOd0FGSGHhRr5ikf41y54dhc14WehLxd2f1pud7pyI2NFRiqmrTyzlMjckz6XnRq/eevIPf
MJUDWyAsljn5/glvhcBBJBJ8pnOTGEYx+f46ug64oj6GaEPAjUhS/0AUWyi2wwzmypFqpYJ9qPIx
UD2jw5+s4lhucghsJCNUyBnApfMliaD4uooncn4XNYz7uwLlzxKDTY5ChNySfevIRNCt1lzpaW1O
OcPY2pRMyl8vlHoSwB/d3fYDai/NvCoZQkS1vsKIwWOJHj2gAJeLlPFkf7bgYctZhJ1Zzz3gwpBE
6aDaTr0eDyewO4wk7vX9sBlx3qs8h3Jrim+iX/leSGKVZyzE6LEjedkI5vlS7FAecOzkuuGlPklx
DV30M2dBHY4wMKnFJ1pPg9rlVYWMYqErKv7LPowAIk/fe4i290DKWYxNQUGHkviuDEtF8YUgC2l+
nX14kw1OIsq/1Snghs8tvlpy/XQeVSCrX3t83FJQlFrQJrtTqM4zw00N7BL/M1ofJuP9SPQXnhLw
NHMoiez+fkR/LjLTF/TvHHVW0YcTB5Vg+mFxptj4ne9fJWaVO7qmWiJQ29MBEoqEKY6Q/mf8j+bi
jjbUXZayhqsejd7c/PCtQ0nCyxbhaRIxog5UkpdbTb4qDAZw/vNKyt6ckx4kgj4nkFb09+qexs5P
CGS8O/3CFAtcPQld3a3vEcOET+qyW84IhjTPZIhx6vRJXS4K7BC9WmN31VVTz+DhcQiUqCsdF95O
5EKiCPHlNYujJpaoYsUPUyeWuNNqljWB/MbGyOZhMp7WdyEMStV2r6yorDNMPlB9M15N6zm9F0kM
S+YOWhm8VMPB1FNOYNZ1iQKF3JhSUWmXn4vSRGpRrTRCDh1hipqqxfGZknESuEHc66ylYR16cDCX
6R0VEVoQbo1/vAl7MU5tXaRW5GIUXDzruc4w2P/TSd6+Yygqb3IWtQzobcXvFA/fe8Xj74YTNk0q
nt58CpS2KsK4+Z4DMeVqarPC02oPZmS7m5WGlNffjXV4yzUHD5uciLyHjPGPY/Bvkq48WeDWDFUu
fwu5fo3O1va8gX2B/TdHNLzf9jW0f6l8AqLZ2Hge/Blvy6ZNfUWFyIQb2CcMUq+0xCxG/arGIPQE
mDYdBrf0wAOZYPC3xIxHVOSBq2cxhTTf9xWNx0uyPT738KONUViPLdK4N0STsP210XIoAECN3hDR
jZ1WuH7zwX7N8PjdUGZKoVGoEW2RbGHdw/w9Zzday5gIwQwVglO1/pg4uX8hZC18gB4mw2lCkMOz
mmEIZeD+QWxObPo0Fv/rJhMSGk9OrZGtGHk2Tw5I9WauE2DBnl/O8RyF6nvQnGFwn0ZSEh4cNiNZ
trNY12fh+xnTq6/4f+OutulpwNT5L02mLEs1ltMO4ncmfaSf6vZgzsRAkOEpdtpEm6rYi/yLTGoF
AzE+eVTf0ow+uJV4vZdUt7GeZedzkEGDk4Fm3CFMQ+9N18XWOawcFOcyfKwI96abqKl+sGPevAuz
GrieZOl/GVCAFw5k0vek/bgQ99NdhIah/66pzBd7hrHhkKCK3UWLhv9aR8GiEAWh1f+4dmluV3PE
rHAQKXpUgSDdDrF9GXLWm394/aBG+H4sq+g5BmQWg7gzB1zGWAzYNN0n2KC2Yt24yIwXlip1Lx3i
OF+6w2oXsNyxDjYTexELYTGJ0BqB3Y99ks39ZtP3nYF10vDRlpyNLGi2K2tLnswvVJBL5qiv3yZx
DQzPrhSDDsa3xHCeDTgYm3FDCnm6ZWqThMPRgkvE2PvQ65ZzLn6UkTlRRjELoirqufa14Hu6jpPL
orVK7cKKWmQk+bXokrRfqsbqPvd2jHomdwJrtd0y2wjefppWh8c6c2nufsZZhMdIabtjWym49Zez
pfu0v0VyFlT+XF+cg0CmqT9POfWvOM5KbSK+HyG/Eds1UAP1BH0K6io6VB8T/I95EQXNEmvVNOWZ
2ijTlqbc7Jaq3XxssFFR+H0BuzCPaOy5qx3pOaQSplXXLiCT0YrPLCqTKGigVbv32cCYCgzzvwaw
ebnF73b9CHxc8fi/Bvhy03V6ThCeD1JWeQ5WfuHPI3q9aABNQYDLn1EhuaFDqHDqTPI+Fyzi5USt
8+Q9EB/JG4K57TQ/lA531l9k/VAV82MXV9bUE+6gvCoPoUpX1EYgD+22iV4+3YC9RYgmC/EetCpB
x848vFWlmVKfiUIM3qoJDCUKHlSndrFC+s4t6s6QKlwsNXOLXHLan1QsRLmgpTwaF0YD5SgkKILS
XZL2ZpcfjzQ/L2yiJCdysI9JJdJTO/pXGS1/Ym7lC/JeannA95bEcT5CqvmN9hi3QkL4uO10EeFJ
Rp3hUFeCKMESFEpBeAMftgX7lOHQii4uT2QfQIACNi06Q9iYklpEHlgcbcptbFev7elp9EUU/ICM
mAG2v7fjJeWVCPNNcLboQiO/0JZPKOv1fbQWgDfaS1vc2zGPkO46GJkaFu6YjEiwk1QXdVu7YQmx
4E8ZnfGvlgB0C8eHepbDAXK1zc0hLNIMoeY2R4k8DjI9FwGCxDYiwOEZVLvZu7x2p2u3SDd28eir
R0mXbtSyXnP2b2U0QyxiFIE6ecjKL4VqcFP7G+p0Rr75cFhSK9RgTtAyoKJSUshTTLhC5xOXwluw
JbkUjEHm7ke6GIbhKUanGVenauRaD1kYqPfeO3TE53Z7jHONPlWQeHFurhBYLkXCli7ADkdtECT7
WxiKRyNn30dLMRg6FNp3q6QkOAAoiTRcz5sFSk8iOtfZf+CJAXgUIxxq9GTXNq+iHX1+u6lNnUd6
8uoSolpHJ7x9HwkuT9qypUjBGmNnxTOflDQt2JxUkvqaN+qnGGNc5GECDhGhoFok3IUVp1B829Uc
4B14RRPYc03SyyliY3ozBodPkZ5UUzUB2briCAoZtWto2f7yGdrD9S0vCxya4odo2nUbq8R1YTb7
bDmtMrMJLC+6Vcgp4fGkTosmPDdWCtFxSIuuRmRUoEi/y3MwcrUn3ZdtSGqCFjJMSKoQ9IzguNx/
Q3YLoPVam13+ME15OwOYkiiMVdv8+6/j4Glq55CwhrkKE+gEaWHfz7fvpkQSghwwZ87k039Gz9tv
fGLE1hwU6xKQYg+s0ubafap3g7uSGV5CKsrc0XWo0yFvce9CHG806MOpyw/CY95qPn8j+5Zk3hEd
CQ50yM8dWECvT/jPo3XUQbfhk1Q/Xl1zBZWifGkAzXp26ZBLsB7CRQQQQCcX1xcPgAjzK4NtpoPZ
IH3dqa38ONBgzocMHyQXjtqLyH+FEM45Qp2u4PO1oU9xgO09ribXpe2CK7VUe8ecYTLwEJXn1Z0V
YfK8Je12S+nnFxhVUkG1IL78uJ9e3wGKkMKxEnCfg+fZMchqLiBvTcAOUV2EFExFTL6+gmk5YwbF
c7hAPJJ9r3SYV5V5Ab7lt106kjmDqQ1v21j7lhXVheudprPajIDS9Y6RE3yeL/QYvskUCyE8KPld
7bFYvcV+NlrPqeT4fvC/XBhpd35cbEOhfnOrDiyJJ5d9TSdfBVstsaVTUq0jzucHGq3dTwnhbX/j
WYeRQk7hwkqVw2zHdl2WVIo7wiCaDHEio+FGI+DjOkfyKt84FoKDSi/S0+eUc4ZPZWBdGCTT8tfc
j+RgmjYI3JTr1BASN8fKRcaP44yGeCCtrD6QBN7kbWfqMO/KQrbQk7kcaJKGxQQiQ4GKa+vYmK6x
/tpqUb9DXhu/U53BNiCf3T2ukRlfI+P4gUbqebK+oikIcRhyQ0FQLVt9NEVLSeJe/B9YEZx533LY
sMk+/04Xe1u98PCl5i6akzqbVM0qVGhP6VmYU4XPtXjYd4W3n29bnb76YygUU/KteAWsCc7Lhv+T
0r6syxxop7DRUqlGCz/4cNVQkW2ZY4LpbnzN9+SFDHrxJq8xOMH2IxvqhrWww9QqUBfBitAEWkjm
N/uuiLPUKgag+0ac4vZrtJOAZ02To+NORPCr79v5NzSstb6fMEuUyeyENVecckiAR/2bMtuOXd4V
LC1IeZrBSaF4lo+05i/XNOClnylc3VBXs6o0vuyE9RXV1OsF/KdTJhLZtgTHCpZcRriBQBZMGB4I
85/R3XKZL1qFXCjtrJDRwdkt5NrlLzcruQm2slmFR0wDQdiyZkxAIZCVJWunojZO3GhLa8RStC8J
+TvQtALvrqFWzhyviqDdwQUOvZeorVGPGTw7vCvobWHF7P0NTBuEFfeFiPe4IJNpZTIIYfKXDm5k
/M9aJxtJugGg7CKRjKWfhxXo/0yGaKArfjWW4m5pixGymVB5eaWCmWzeLxeXNyIhKbPhLWGLEYRK
JGCC9USZPoorZy4RXobdAPCMnPrVVPpWxaSJZoBNMnvS2WwvY5uQRA9oXT7Z0xZvtmIz72BJ5V9B
zPT1eF8yKJwEwGeF3UWIaZPrL00jRUuT4OvoaC7u1gjfAnBn4uRA0VC3TB7gsnmo73F1Rlt1uKgl
xdQpxAlopRygDfSC87KHpXL5IsAOJaTX1v7xw3Sa/Av/pH1MIAVN418rykvErtOJAXSQtv5gRjzs
TpedQTFJb52ucqksrY65XGqeWdimLSxYy6I33JEAS67hzKShzOyGgTIROGEa+YWFJT6hi5wBpvuJ
pTzQnb2HXlw66dB2NjhxYfE1fPmhaoQgk+d482ZvpoxnC+cKzzp3xpyHkt78hjxDKHUgwsosfY05
0wd0cKVekQ/bnRdacfOhgP2YtQW40j8LyNPeyJDv9+GSQ8xUHXKGcFTfKs+QZkzBovbfm//FkR5x
+MK5THE52LV0AGLiqZfK24cpkkJIzUG9OfLIOMcRPF7QrNRhC4noAlYtOZuU579YZ9cdsfK6z7qA
QyD1iYquNGUwxt6TrH6JppJVdIxH23OYNcYmBcA7L40BQPzfyfl/K+Of6aJc5zBBe1unD4P7MRsn
FafF3XNxhvePJ2xVH5oieRhO/E0MHNue+/SWB27La0qlxA6q3w84DYlU9Du32n9BZ0yDUnZKTlcL
mJBeDWnvXWcJW4CMGaBUXiqJhXNamtOTkyBPaeEcd9mEAeNqCzzATaz7q/rNEghLbPEcwdyAu3Je
Mu2/eiM8hSdOKaEMlCPavHwPVmC001h6p/q1M4JPySl7k7Mgo+M0UnyulMZMtjSTNnBwv2fnKqqD
gi2FPY0d1n0rEueS2vcZX+ZhxXDRURErBxO8sDOAK5E8Y31JrpEJIHMru8eiJZxRv/QlmPUBAnOi
gBt9mft7scj8ycz/tVLwDZ3CLA6g1saZqV0YZRAw0oE+fHrlNNGLEvcCgzDWJCpjuJfv3Ko+mfT5
nwy4m+U3A/FKS3m5jOHcu3LAMhaYQUkv9PurdF9jyciZIcIJDwOd+WzxaBdhHa3INGdgDqkuUaJS
UHrZWGnEkgGRVQSoBXNyugLvHGBPIZ1DH2HFSmjwr60QMYubOYHI3/PCQ+thFv/xXMxPfmIwBEBs
1+FMyUf3riQOpkrWK3n3mHdM/q9HQGJzlfYhb2JryGLXWNDHNvV/pkDZcxqJrO9+06jf9xRRsXXt
kKcGGMaKYdIs6SxJUzxwdWRTiTE7y73OXj/qalgzCg0eT90VqKIfeVDUnviqQKznnLFuFqBRmtyz
DnZrlw1ByOdXPDboy+Xp0onjH4Lf6mqgUG/2q+fo+JvCdXBb8bKQ+B9uLv+cpNllGT9MFt4WYGbm
YcS7PCJnJXEidr7rDJws+X3tZYe7kdWtuHYeF9h3AC1+V04v535na0V8btuZXTP9mRVI7R9GUjHK
OFtHKPNec4sMAt5qvClDSrixkdksNF6aTkdmLaQ52OyUrCX81h0oHUahPtiNdSTQu+c/mcOeNVzN
fCBtVgrqCkNWbq+opAJyn82B8eFj4eKAQQRngubyAFRSyIl+yf+LsCgBRM1F2ai4mpSCCGGCJ4PA
iY+3egSUd9MdUp/MsKqKW9McDrPMheRhT9r8LdCmwlIi/niZmg8haNsSEG0ipExdh0cYxv6FHsMa
BppYvecJurh5+Cww1tS8dtFD6LRWBXQvggVbLNuZSKjh15ewVOGQ6/jLk+wmya0qGpcAU1C5TrSn
cFZK2k+Y1WqCJdGfQLRBKLXWcfPGb+bXPSq9fVQF1+HEA8h9VZxpW3hamOOw32GxxcqQVI51ZKU9
p6YNbaamnJDl6vtaknKWWQezjV7aW45pkKLk1lvDZfc+Ej6clwFRuuIAsdOQWnGZs8HVQe9FHdQO
GHeD5RjHQ8gs95xj7I2BQrUHrq6scoEPcay/7dEfloCwnnOPiVnnGwJ5X5qH40ot/maizPdl9Yin
DmG88UIubCNGVefSAwJ7wJNAEsCSJg1wdmDrLtU6zt2cb+v4tnEArwzvPDmE+/jJNZqrorHUZ52N
OQKq1qNWHK+rY792nO8uUdMFFIvgh2pw42ljcggdFoaHjcOvnFd1sedxtjPxPU7NWkThtno1Vbtl
wSolu2v0xqENee5IfX1aO9QU+NhBolaAVYCwVMX+c/9wpsxO1WFUjQwAiHYQdNtlfd6o2GHtMctN
cdMtxVCAHJxoYzP/e8VfEQvhSUfFdPkpUAbLtRwHYt/ZstXz+kP1i4sf644i9QtXq1aT0lryxUX2
Ql89A7/2S5nZ7tNl4LrbHf6gG66OIdAwbBN3fOwUtPUMccW6AnOi/MLiIl/NfM7GUCdtHPooElU7
tt74t5ypdzuDSunYtNtWXD9wybX1uu4h/fhEtQ98eQ1U4rHzqqTCyrTv7orLcbZOO4T6N38FRKKm
TnIIKCczBjEanHGafl6sQymR335PhcDsncJ5lld+ly27ryMxF4Umnd0wrPnrR43vVaz1ACbuVdTe
jR/FESh/cHIsWCTmAq8G9AQ9rU8ye70QF1H6BdBDBAk0c/fLbyODF/avU76ZZ/FwPCzCPbss6tx+
LG/52Y1l+Q6DuhEY9ZxRQ/5pEEbh5udFxA4BljlIWTXQDyaV4ufCVYTOmQix586CaEhaqZJJJpD7
p2w6zMsv6oyYXT8xSVmDlGokc0MKdV02G8DP5MkZyJg1sdJ6yTW//GaPv8Rx7gGUFKHRZCKvjxfb
7CHMrGGkSbf35bYeL8AL+2M6r5xZFDEghXm+8djQvIpZoxfU4Ag9IikA0fGmVjYT0iVHRD5/UrVB
isy6jDGevOfA8Ldew6nQ+K43G1PA3JX6rb24Oni2qhCpXZlBlVHZNEa7+1KEtQJBy+/WxeZf08nd
AXUGiVhcm5wMzVPsk0HTk1dF2GyNMUKbzRbUNZAwnnFxcDmFhlzFOyP1lGKdpqXxV6LokyYBkuky
00VG9bHw9yQGCk8pVKKq6/7jA6wfbazTyLuGXTCTVbUfj9RE/yBIU3LruapYt/FvA37Oj8DYFX22
v59fJQNB3SqgEfK+rITX2cmgG3pKTjU6PKpfHelYqcqZcYcGco0ZN3EB7XsiekgqIKpGBUp/bpew
8bnYDQwkOwP+oZA7kzcQ3MfNxBSmn2m8/W4sh7xH6TlPfE8P/LLjY7x1tIvWSXoA8sK7LXMA4+YM
ZNgyNC6DSyAxm7MbU7ht3R8WQxLz9cqBQoqt+kih/VfLYBZTKf1xtQK3JA6lgHpG0a4yFGk5U2V4
gncGaOMM2f0e4Jgiv+ZarS6vQe+g5Pbfa+rVUC53Zd8DFaiDsmdx8z9/LB16Ao+lr1Dy8wLkcy4M
TckfDk22ACYDo/GYtE4q34/XHkBtcmsv3eCKYBU5wEsf701UsV9p3MN/pWidIFAHf5Ha7ogMwmRi
RZjg1mlkFBlGWQI1HkvxKQVIk6CASAiBSVDI05PVS8CATnEeWWrlYhnhEyyQF7HVjOwxF+8UCsrK
mmrSUYwXKt7bInTZvu2/22OjqCWMqyBN1ReABTSapWd5Lg/pL80oaZE4qKk273JBOCdsF2QK7ePj
M2zFrk1im+07DRjGwDgJeLFzJ7dt+fEgY2prU9MtS5Kbmz+gwXdidrGymKgEJZMAIWnrBGv97XiT
CedCMKg1MUFdgywJWxJEYy96Ie0WRc+4bI1smcpIjNyIn2TldHITzntH3xNcSaMi879SVKUfIk//
DQb+GS2hwQI1Dw/aPzu2JXKYT2sLYf/8RZTBfN4aZB3z8wn00d+2Youyaqw9TsCCRuXofA2RElLV
7Mq2TH5xWvGGL7mrCwT9m96S48cnTZiUWQ4xm9RwMlnbwo7otlfUVrvY1cHKTncxGgf+C7RlxDmg
CdAay9KU95hiAXee7dlxef1HgfNoa+NYiR2Zoi0jDtnbxXF2aevlTcixkdgX3xNsZuz6gVU9p2OX
m8NplHLiQp5GiBnc4Ue9yuhoUCuZgFnK0PNQ3Mj/Xkjm1gEWp7GmITu0QQU86PyNr0a3YtXoXNsb
/zXJSDYfrC26+wHb5urG/rXG5oBIjXBc3cUkN9RPmHhLPt0lkfG3EsnfKuux8NXR16Np5HS7M2LV
UomNRkZ9aarcEs09Z3gDFF3jkZKba2eHfXQi+2Psvrqc/MiR4Hjor7aOqkD6lCLY7SG0tm6fjAkd
+Z2m2g4DsIFMmuFAbKKZ22JOh6UbRVBM/pEj0K3JLkf5MK2DqgerCZviB/1oNdXW/RYosTU6D1pN
vjvfTYMOQen5lL6iztNv3bDwRwtjad+PqKpPpjEsX3t7itsKcvImEICbmXEU3/D2soHNb9mlOG/O
R0olAV0zL1/7CmB8nTPsKpEzSTgCP74TLjanaPirxke9CVWLu4bDTvRCB4WBXI/Be4/pzyaKviGP
dsPofi1hTI1MGtWRJQ8HN/hBxqPuZ9PkhyBkUHboy8XGVqSFI9EpVklSGcyqPDzUnJ6Uc7PBOu4E
pBeTUNCUjHM7qYAOTrcbzkWVgRyr1b45EGLB+CVQBBNpmOlImN/u6fkvIn1Z7cEY6o67mBeLKPCJ
XHkblJafD3RTZz+4uALnnVkWIBdwTiuz2Q1IUOBkFYwLMFsZbs3mzDOba97uefR1Df88cFOT/v7x
+cheirQkCPg87aBOXwbG90LDK8WETmHvTBrWiVtc4SJqVUSDVe+acwbenfCp4j+WGgTwD5FN5nhX
NtnLEjXiwWR/gXL0evyJeMiAaHHodvgVt35iNNwGi4dIK8ycL7Iv3+zyyhnqdKIZpmi15aEyLAMG
zx/6Ep4C4Jeyxr6sKpjLyl/bkuj1cAgGC3zYbwESF9ujSnHrABfu079Kv7ZDGsny2aRE4Ew61R09
CufZ+Fg45io2+FFHSxvR9Ym0DlhG5Y2eXGlN0KimpKHXLNHjAxJ/tn+m9v4Y8DSRN22EMvvOSLCO
izo8bmDJeUCtkpnYOmu9lMg0dG9AB4eApmfRAUdPGmdri1jNO9kdJQQU13irD5ETDjVQtRA93xbR
Fyw/q/GTO4drMeIpc+OtmNt3ikVlFfIBbiK1SI5j0KdEyTVUTVhuNRgv0odLKI7gzbw8iXRb+C0c
l2jE4bO8kWjqvnNI79mnOdVRFLgWglTWvGvIAoB6wsxxutlPr73+/RU0BPt55wnrp6J5+CokNf5E
PtZRWO1Fejlorywhj6CUicZwvT+EEZdZYkfU1Nj/R6R1hx0KY6DN4PKTTf1qZ5KkLc7E/aiZS8h8
TZGrXOd+5Jzsx4oQYJ4B46t22oiuR2WvzahZH4waH+RIqRuMN5D/tcRhfEaYhFopvOOhqzqbZ5Db
v1lQlGhCTDF0vMBvCYkutAbJKs3RNXJj11ryGTmyCtWkkqa9br3VvJWrbhpQQv05qQ9BgRADuMn0
eGLd1oKIcPWCDTeCwHuDwvorbLZOJNG9i1g6L6fzVhXzjl+tYwpEf2HnUfmCCi7JTSjjx9CNL5bY
+pu3d5sDcToaNNDouv/CeHowu60Bk0OnBH6PS64Y6kxBDwuV9AkkLoWFDnsH34ND6QxQRwUutSca
R6WbBP9RFaJvxRfhuwa3yJyXuiOtisdHdr7BHRmCzSeLirXNnzMHcM/zRzeSkgPulqi9ifS1mo7q
LDR7upSR4QB1IOOcqeqH7ZtbB7pTtoYhHwqszjVSLcC6a6a4I8UIQSVr4qqtUMdzBES6Fov/kroX
l144vL9Bp/rg7tnqCiX7jXxw/RKprRSzRLMBhD1uhipuwCNo7V0uFTr3sO02WsOCakmxxkQXi4xV
G9wfZrfCKG/Fo8Ejvac+slO0mNaOxY/NYi9N+kGHMI1N3uhp1llbymQbjjtnd8KwdRhNrtlkp3QF
IB4VHmb5qENWEohn2P0pntMbXJhIpSmsZYXdf7yMuYCZeI/G2S+juU8q3dtR3FbDVALWdX1Kzpc0
uWwjF7PWIIOHrlEtfRbwj5IInpAE980mG2qZFgkIhd4z5Zz/al/J+g5zEaLrvMSP9kwSPIwCgzNy
JyZzgV7xrCjDV4FqBZ/mPDUTQQUr9SOOPYhy48M9QKWPfc0YpM5hFZwftfIJW+kDK0/T2pkSLKNR
khOz5k13S0M6vUDQzdOv5fAlKa4GUX/lu7M4w3MWcpqeVqPHxdPiD00LAw3ZEi+M0576NxLR9mmx
YmGphyo+KIFLej4Ol1hTmqnCsq5jCixBKFZHiZYJ0A9HN7nVcyjyq/Ac2bHzjhx1BVkTOMLAkndv
TLYXLcYOOve71ZjpO9+u+KVzsQshi79VfU47c24xYmDuu6UAvycz/64//zJQDGlT2mVipAZIJCIC
TSFu1gwoOkiV5d2o/01i9TX3oWmzXpVr6UxhRlRZmG5QfLggesgzMLykyAB/Qw4F0myWqPMncGFf
F9kFDC4c44j3rpA9h54y5b52Wk0jJxOSafVzUU/mbNqI5jNxDxJp2cdM4KbDP3nFtd6rhMXZNHvH
hJ+qKFD8DiRxYKGyDXEwU8D6z4T168jaNNOmz4mvh+tlsIe4LvNINuHL+htVpgLrGZXOwtx1dqe0
1JA8h8WtTSOtbvx36SmzrPIk8+aQUhueShsdYYwcCzdFh/XlGgRp/wkriU3zkHRv+YnRPz40z6Zd
REoOPWVIUbBKHZFlPdpEHd8d8fcK77JMbTe9EK86B8tM0G2dckC4+u1uMw/uX8EUubbWwXSeJrqQ
U2RYwggVC20PDKkSBKsLJVQSxrr3dZ0+o/BuKQqgSCuSkpr8+psrEQeXnaffjGpzBWN2hUS2pz6z
mQfSKSr8M0W7mxUwS6RR7aUClTtKEC3RlTr8IifjN3jTG/YLxWcfHlACjXQ8S8OupNzGJlZ+OgGH
1y1BPd3+R56tpdFSp8hxBAQKDOTVhgFSqc61tTCTCH13V6vRoXLvqkcbU4EjBwEkVDGz1bhebRXn
vqSvGana1zMSkARtlJkxy+c4QGHT4wTp3YobDSDiVHxDpCNiD9151xK2i9YaOh5dyS55a3Z3izDR
beWgD/PEIeRXSRYdb/8L/QruVC7iiZR5L3Dh0bOdBnyoZS9rS/tThUukzLQ+168NDdfZqw5TLwh8
mQ+jqNxaJyrB/YJg23+d5PHS5eysvldsYHf6iJA36whlnNKRfULpN1ufegKOtumylEEFYbz2T1ie
atRHMYaxUlNklhliYiqjzyAVcO8Fc76gcvuPXIvl9xm79TScj19+NnP3NXE8ijFNkV5oP2lAkugD
qZjcFfi6B2pDjT0dlvogiI9p8qcyXCW3LIfAyTxb6rkSfieA5reEc2jhgq6uj6DBetmIRckFAMmD
tabcEaLKDu1vj3aVo8mClQxJSjC9LrJApcjZj5SvlCesfUpZdptP06uX+hg0s/+xVpLLNtkE7Tym
3J12axU5ENaJm/HL6BL71tPAfEXwS5D8fYbgubg4OStpiXRGT9bsbfkMuXuVatzSMGUGx8jrCDKO
F/J/VhDaOtthctx/tUfMR8Q9/fTZK2nuG6ufVS5BH5ylDQtLn9F2FUyjpbzZsWmLAKB+qCQhWKs5
TJVyJvnAGfR1q6yh5eh7latu7NUL7wosuin5PHYFfk/eAx+/QwYRjvQE7rYmHR/zLgW0V5pGNwea
WyKJCyIcw1iO+UkNdicvvADRsEP9Q9agJBg7JNH5U1X/kLJniU2LngiAX83EY96XfvbIDMm/So4q
JI6yKw+yr7YsDQjxaIHfRLMp6b1yhfOJNEWmz/xl7tRedLZ+t2YgpuwUqeQ5+3MCGyzOp5rJG2rb
/6rzUy8zwmKj6Ck81UAENERE5qOEY6HIO+nuWVOlbaTroZCUgE5/B23EgBIlpMEEwQkOX+oftrVu
/rMZ3dQMdXzb+DPEyOgMZ4H5ZW25Ao3Mw1R5Hm1hv7RenDq0kbJtFd0r4Uw0Vx72EIEeAA0WvU2h
e7T+dBuAQlCjuqFntmrLukVd7RD6NjLm/LopdbnYLhp9SiyhePZXwX8OaDtxCEjHKWSe2vkF6TAB
hy/1QB08QlyV3BOAn8R9/LN6A8fDmXUSxLGAUnYF99349tLltPEYFCSxOSmYytGpEpOiQdRL5v6E
RloheoHISZT2/wjmy+MH1FdN6ydbPHh+0cF/s1hB3koaOYvOInXBDnoPjGkNiNt+xp7A2ZXNPF16
esAZMBmf4SvikrDb0so1+YxVvPOq36yPEHQJU/TemoIgFKsR1ofDMgDahNYMCVf6r09gYYVXywyl
HGDSXJQZpu2t/+NFTHHMEZhGVW/kvLBEDEsqlRRxRi6iFg5TILVieaAdRzX57CbRIWEP5ZPjqGGx
zU1DKIQCnsGKalRlbzENe8YMED2h4L73nPsalWy20rDKHnyb2Y24nkZ3+tapNROPGDWDA22jEBsE
vZyFKC7i4akgBjxujkURDCKN9ws1F8fxGlUGCMz1P5eRb3IKw0O/Wdt5qHMiy8HC/1zd5fJLCWeo
JABh3L7Nj3FYP0DtvFbi3o4WmUICFQMIJ7yYqHkvTrwgSVNf50hJtlywr1VcglDXMYQDR4kwQQ08
jY4PCHNaZ49u6i16aP0qSNPq4uq2+PVkiWcHns/vuyjG6gB10ezAW3mR1C87Xv2rtLNp7K+GBkCd
pTeY5+lXLJFK6H9hC8HiI6uren5dHlQCb9w6rID1ahHOUCWw2yzTweEaka4LLNt6Z4Y3De6c3K69
4Cx/ofynVAk8EMqA2dZZ32ICEXjf3aVbIq/asmVe5cf6xJa8KgtxApVd4UsWZab9kpYPFlClzb+1
KR468YTjAXU+cqe2j1bTh6uOvFMDSyhLEI+sQuTGvhIspvaYpPhf/ucJCxE22J5sZAHuol9WW1tN
qx923aB5s+d335H8DzMGsF5yOZwlRLkBjH4YCL5bB8wlowDczBi8C/A7ISQzHnrbrvxeLpyluZzp
/c9mX6kU8vNsUNzSB+P1BqKE/EzJmHe4+R0ybYmAS+3yvHa8q0PnEcNU/AfsA701S3RNC5T6GCZy
zFqTWN8bvZ3euYnSLJnUavAX5ZGro/Zj9MC2+Vna1HLguh5caJCkGZkg0eGaFHdMd3vSAC81ncf/
F1Po/XRGMcmQ/+QZNA/qjq4MPSgSFQSSD22AMbelXSySeRkkeLex0D7SlAUoI1omUVVIXLlzYwRn
yCUle/xBx56chPbrpqf0cHBvDA0BnEAb5WssoML0sOw/cSXjwarmF4QzA5KmMIIlQahG98zMLOXH
5HvwOzUdUyH+cU8sCtr+yx1Qez+mHi9/fFIk3csQN2C6eQzd1oGZLEcff/gACj9QXc5hlng+RGIK
lripSHM+TB4yqag6rTSpsfEZ0e9VQb0lRNW78Bh7bHzqDWeFJjKIA2WwHfTx+0Rqq3zIALi2X8PG
/DeUu/OdQCg+tjgHpHTaOc8/BlewqgBvTi+rAYiw0PhEfaJg3iL6TTMp0JYPcyOHcYSxO+suZPy1
gSI9x+XhT3dQQNiEd5aAigwqb1E8yXs0Z2hRJ67UP7spHrBLcAdWv8U1JGkeQggAM8wvNLo3BKbI
xDnq4yzzgNQjlSuUNM0WOvEK2EkMcgGZ5DvwbxonVfjumpJ0JyralSgMpi4uoMablILLlxNb+EAv
8vcGoh40HWtKzYoFlyG33P8++sZLiAlQeTkUvPd79MhGE8FuDHb0q21Y/pnGUZ6c1SC9qTYWFmCt
4G1SM7QqAMdkJe//fCIvf0YnqeS8/BZVZteniXNGcuLg18prYD+z7IQjwdQPIv/lNGi/eg80p4eK
lsyC5RZZ0YD0m7J1LKGmPDpYvuP8stX4+DjdlnKOHM/Ui/dgifVcFIIGJYeeVdwPqutWUiLG5Xqb
urupoXV1lbuIRTJA+gCarkJdzYbRMaEWN6lkktIdNlvLmnrNGbgRIQeqrbA8vvCHU12zI3JaBgh5
/SrOZpp0WS9RrYYisI6VTxDvQVEynUx3glB/c6rxenTgnPV/IcYGKlLqaBu5/WSciSfhyOH6wzOL
2ojcFqZ74LmGE9CLplzJdoBJ1MxgPAFC+ftX1EAZnXJ2p0LSDbHRYloQ3m5+GrF1g4aDClMf6cCc
YpBe+fZoRPCp1b+9y0P+eBvbkK/PYCJi3jMGsR3njzzrRiJDRxR/XrgMTIvGifd8ehvue61a2xDM
YUXzj1w1J0V9sP7sB4XJV3+/D2WzgyCh3XNrt4igvMpPC4sNyYqfuf5azWjti5NkDFVLEyn/PDgO
x3kLA+v5Ua7rmv5+y0ws/NPishune8pfMyhhwtgowQfCiLQ8uxisIfIB/XoJJqTwE2w4tZsH8gP7
jJ+VCtRX8+bR2r9MgFFaOy6GWCjWd7lKx8YLpZcWY6vW4cJQfcMr6SXT2oYkjB2p6NztHgKt6dgy
Cu8kNRDBjwTa+voNANlXC3WqvqRjYsqFfrJIq5n8/+zddHkVzchHRWs7k2mkr+0fdA4kfb3ZSuY1
FIGRtQ0eBWpMlOY0i+3+it0hEuVq+mjvmSI0otwLsFIq5dkp9gXBzXPiGx46RBvnSWMyLLZNYzoG
O5nepdhDVb8kQDOo0b6ueWgvMNNtfH1tx9f1DBI74yEHsLoPje5yfL2XGWKFevFTPmu1eYjrBJP2
sLI9EqljA3Uf28YqDUrml7RNpqUgt1k/pkSDxQoDo7MpgsBmfOA1Pm25FIANzmj4C3dXmN5V2Dlj
q3MgvM//f4EgChZ+O8QR6QFDtEuSXUIlXDjqffI2oxTVlbFlBOCW4SuLr5FxtiviPqR/Y5DoAmxx
uwzsOQ2VqZueQMDoqw5ZNJ49CSn/Am1mgJ89aAoUBZ6nNygdYxAI7pR6lB2UN/mI6JyCT7uXymHo
jeMUE/8JtQZKPDPaxW+UWwFNw+GDMCvUFE1vUp5XiynTxxkzP3/sqMXKhJWM/duCqcwFuhZhwSsZ
TrHC4QPya8nIVMdcP+Iz1Nzqi/YrEQg+U33wQnRoFpkQgMdOdgoLzRWUCAZZP/RLHFtuyikGdwnE
rwwtKQ654RIvoCGuJNRpPjEf7BiIZtgNFgt7nQa19ikTxMAdjCrLm8kMIqoy8E1KSyXDo8xvmfsn
Nv2W1ORxUgjlrktiFmJ7lK1uogcpzAQ+bfh0mAg+0VV4r5UvhR1iPEJYYNxCSVnBQANfh+113xNi
1R1bh3zMnjcJgzBw1gnef4c1BejjfZKOZtIC4NimnZGnAVh4qLQVrMytgfaWzJe7LVbleRxLt9+I
pRcOycbYpTnox9xyCLIXMt7WZO1NhUeqfeMboCQJ1aj8MN6LpYtz/dT7jkJaicwys+sM7/i0siAK
FoWu5pcXcxxJX2VOtPeHEwp5j1SXoVdubumhG00W8HVMv4jtAEav4BQfkp1moC8beao4YlVtK54I
JHSCzJwrJbkOGq5L+p7dwYQHWcOMKyRXZFQ/bTDEEEX+9hsS65iH2pgbcrc+4QhZLj61ocxrY2P8
SsCB94toSckP6AuQmp0Y3xVp1qst+15eiqk6rjdQ24LDbcQVx64VLQEpXdlhmGzRoP5V6vs6m/0V
yxzn0++ipt/g9Qkp1AyENXZxRa/qAw+bbuqNAXQ5yf9AWFqT2x65vvizhZQvRVZ3c2ug+PZCnIel
6+289M9HWDw7nPKFNR7KhkcZpBO8q9t6sTjGeox8JQ1btzJrEMU1iLaoyZbXC2ouVTfLWbPifrQ7
ssS8B3TmdGmnDQZV2dtKLIKVzs8QxhlYGtPpt2PDUieu0Rq7qIXvXcUG6+z0EwzUkfZFqutmd3Nn
xiVh98IN4ohjBScNx9XfMo1M8fcmXMd3qMwHNoooJiXcXH9wX5fR05zQmshM+kMbppQtIkJwLHAp
tHCOML+HUbqPLTPzv/EVkJgB3Ah03oqcpUCiAjVJCW1OsP9U3tKuN5iil3lhH1h1IiA6W2AtxdgH
DDXuhxs67ZHXeM0nRqO+9xTwxR//1kODiF7uOAiTE2KIPXtzghIW5aYJ1mz6UxJFSD+AAoncs3LX
UgnzqChksWKrUNNi5XGWqRNhKuGD9B7myOdYma7QlUMoMPslK30ImHtmgrsy+wekxLbGmgZHWDcg
R/NShelLrEu4O4ORNYY6cMHLGrIZzYkBL5JkPhbAH6E1mBP/p+knZwzyOa+fGLsCCnS/dOtMFwUH
8yNhbVzEDGDLTnzewVIbZoFhIERadihE0mODegrl3f7qR2GO94qUndVlYzctcNjXN/l9P4AzwuOR
GOQCxgT8qhbk4QUAf7x+BgBGlY6ZrJcL6B3+W025T2ZV2nDJkUL3L3ZMLkkSvN7vaMOvfyEurVHi
W9XdYPJL6lGQGNOsf8KZhZo5u9l7RdXRIZj+exEXd9R/yxr61kF76+hcRTGuAMkyxIOpsIv6piWF
wLCYNReda+vC/TM7AvkYh0T8XyUDixW8pihFVP8k/3wlAWJjx2d15vzm9kcimKOZgevvir1PzExC
9QXk2bMabfN4huRLe8XjDt75pCjvetXN4kwtqkKUGHIvPQcirY3yGurc7V4YoDtJ/a6C81Rwjfo2
6+QdeEgpyiV/boMeF3IRpVeGQAOQfCf1tyGABqCm5ZuZcNyDnMd5LvDV1eO/nEh9aTIt9xeZZkjz
T4H7hAbQC/sQsPiGyZ55WZ3qnI+NpxQF9i5p8oBOIpIh8KrttCzOsqFLAn75eTtO+Ff3zlZL3hBv
vugL7V6769kGfBkZseJG5cw4aWjOQ6qqqt4oTlRsQjioih0Minwmzwm+gSn60zWMaZsM4drm5Q6O
QGKzo6i4QTWPxrFbJX2owzMi25bKpYjPzAH2qjzwJ0mwXii1fhVq+8t8SkgLWZ2cguO7HMmGMeqd
DztPiXnInPK/r6CfpR5rJT+hZDUnCeKDtB47FywmhBX9OqQPV453RFuc0liphUT+QfWpmOtbP8qz
Ia+Wx6NilTMu25OLjxaD6rPQ8Wt9ALsreKE8Z1MlEL5GsHyigCqbP4DWM5vANSj3zQDHPUPuN3rE
tYsM7aqwRRJqILEe6O/7YT0SxeRmLXajx2Ya/6HJD6/K7WQgYiNVDjkJ6A5F72jWY9IY5cIPLu14
UK7LUKrrZGqJ8Rey6SjuibljWVMR/29VsCrLjpngcp6T/1yS30iFzQGOKfZXLcj6i2akjBBSnJQi
VXcexp8zVXQOC5izhs3nlb4lxk9RvRnSY8oSkDKbekcrQD765/19n7u1ZzTEZoUjnvYxkfSKMVKC
l+Z/3eVJ75j+lHGe1orhYE2mOPq4TKi2hFQHT2Y6HzXkS7Bs/OxWO5Y3Dn3BcSlks8GaAqJxJYKF
WjsjAI+q8rcRU5NFtqNCszAzUHEnvW1/vjwXENTDBONZs9mzTiqKRwrBCdRTk3K61UlykFXAI8Ib
6VQqaQiF1mqiLLRjF2Va2qkEmmDfUeVPgkHo02fA1Fgxck+xkzuhRWBKYexHeC/F8R5l+QQs2s7s
utvoJlYrd3UV5E/LjADXic4ubWuUj1kOR+6EZ0WU2jTuFDYFAAyVss3n91RAEe29b3GCIqZUPmbS
TvA5tjfTZPsTaqTSfEDe+UegHqx26+wimBbLqjrceW89lCGCsqIV06oZP9QytcFel5sWV/6Ev4eb
oKOceLsNV5sqH+nsOaVrjqSkk1tzRmTRhAsssUtzOsmQhTRsREU+/unRyY6bDgJvEz303VcQGpUj
IXB8EEDFqu6hokoX6qFu1469nvwvtSQsRgvzdzI8sm1YvVoIN0CU6XX2NZagUSra9aMA4SioBgD1
MfNUQbfdJzysI7F47M8A28nKGWS7sHAsFJMBwNlTSmD/eurj1+4bF2gTSn41yyEotIrJL5g78870
L1PY9+kFP44ULnw/8C201RBq4tQSQmnNZWDnNI6aicWW2l/eq5LmSv90fwZ2qZyZEiFiZ8CTJLO3
hdUPJ9B4436cTlCbpp+9fzr8XHKoDArS4AtJhvuALNis+xenopS2T4c3SEHqyK3C0e5HIAKr0Ehw
VEZeVbekdfRb0QMTXD8qRYGG7qRUXlKwrXZ7N0DmqYFYPlDY4rnbv4Uh3n0Ac8yTET0GJC0p8KeF
nJppaOCkcWx1SgthCosXHDYCazP2y+D/6fMh6+0PFvgB9sInUE2FErbwggiHaeuoFJfbYZhcdhRy
RFJ3dXX/KvT/ZsV+LMXVgStnITjGf0hrO60sJ3HhrrhBz4gMhYvlXZITczB9ud0fb71WlFvmHppL
YsPatCdY4+ZcPsI8TcVvneTcyAKiW2TyGxWzAd0IoCVoj+CWUXjlJoVS0smGqkOG7+OWDVn8/z8K
9B161x+RMQW3uyGpK/9PWkGtCaMdUyc5n6el+CuFqC4vDwhKPM+dm+bDc9iMJjFeq1nzplXbf7WG
7dVVPcjcVodIhdJASeLeRL0UW/DhdhRcSed3tHGKNJaJasW+CkZ6zCd8AZfzsgOXeY/T6tKxl58c
7jfpNdGa9z1IDpXgMly/QXoE4jityDs8jPK/ele60D2bVr4TMpsGg3wsf2UAqYn/gmLVtIJa8nuV
9qot/zScQlVPxuseHTwQ1Hq0qF2mCrwkOiQk/A7fkMIIHBTRlGI4dtyIWAP1WsDIZgk2huugcqi0
FzHaflX1rvGIl1Mv642Imb1aZRLl/ks+gKbWbRc9NGSVJzwf+pPXDXMNnBU4WjWieN4g93Qus1vD
wy68dyz0n091dY+HxShOkzlNQJWlXWP7Up6xcsXJ9NlYN30N1QmFPWD/rElOQtiLwW+ivMfTfhdc
vx8JxIQ/Djq10R8e2i/8B6ZzlZOZceBJlEAttVHCGLtlwNmJ7l5hDYzH4yM45ldTUlqvjrBacqKI
GVlKia8Sm+EBD3pa3znkaUNAAoaDlidQ/4LQ4Ig71OabYwL/K3zVBDK5crk+6rS4DtDfFi65v4yq
e0xZRaPFHF67XmspHTKaGuOHGvVPBlBvRqKacKFIWuilDUdwtEijj4iixc3fvUeXsPc7XDmE11Yk
i9r3cUN8Wp6I6/sm9khKe72ka2cvl8Fw0LVwa1vP3Gt3ZM3zCHBTAC8+//kZ2s4zELccihYwRRX8
4Sp/XvWcrEmBzGwPBl1JugO8mxa1vsYFu0c5dfAuElz+hMP0ZToj/2wDRHA69NefRFlSuP2z//HM
RT3lSXGAaTjSXoqu40ZEH7v7A9ebNpL0wRy9XJRQsuwUHiOqyf0TojXnMW+CEq5AL7fNz03RoH5n
erRrA6JJjf46a0o7lzIa4CVj7U/jx/OZxwpJnlP+d0p++8TdAIGzU/O8lWONedIuP9fpRSmFbDwQ
NjISWiGYAcfhIisiB4bdc2IyaM9y8a8UZ7yqxZAN9pxcZMrsje0lha44V+uBvKzysHRanou9et1G
Idl4wJpxdWbGhkR5k9v2/UeYayRgzBk9vjJuQg+7ReXN5s54C6ul9GuSKgcC0rDrsXVuCNjoPCVx
W/WyI8dSxN+ZJPgkzaiJgU8Vs77DPvV8mss0nEBpvRdARuR0MIQTMS7sauEp9OF683ElkZittzPm
aJ3fwfERw7JlSp+T/ZxbBtGldWgP1Y26jmRVRBPGhSdhZvHDxxNTgnG1TvfafR6IUGVq5TRGjZfv
qA871Lv2niC3PTBbDeN58Frv5eRtsPa++V6A3DoCo5SBacEq87XMucVTfIt7ky4xngGS88nga7Rk
3mDG9hi2gL0SnMzH2KJp33GJrZLCr6KQfsmSxpPapHSQgWHRjbBfan+b9+p73RTL8VVGXvWHlLLD
LYvxujaeOhowYuuV9pR5fpN9KpxmEkApicGZYsXgoYP5kQCWgNBvaKGwJzxpuGNid0SAFQL/BCuc
l7m/XVNBCKd7ro8ATyUySKpIU6F1oo/KTsYJE65CSIdjNkttKsEodJ2LM3qHtlIKeNtKbPegGmTl
LlGlcaxJMqtNHH6lzwgxifnnbGQosMkH+6N00/+IEvKeZ4zux6fVqBDo2d+MJAwye7TT2tp8WbER
hsrMxcREQ19kB2XT2+tUvbB+pslaSbyhuM7KTIS6n5i6Z0/GdTzJngssV/Rtx1OREY7qNbXE0RiO
1r2t8h4SmcFNNYWVyrhZzcbq9jclUSmNvmR48nfJVLYY6LQgNpHP155ECNW9UAhzdXW1P6eCHAyN
HLUv7V2JrFw9INCYraoXLXtIV4L5FvOZ3bHPAykeWszBE1WHkmemj63qGKhrZh1Bi06p50bwWgi1
HEqUgrCXgy3ppHbg+9YHk+LCQq0GfiQ6/4Hbtkl8Ro5WcN3i/hvd9cgMW6abLsYioy2UnJZvmNgx
4ZUiFi9hBPhqwJBQkaL82sPLDuP5c3+Ph6c4gFk1+w2ZvTJeQeNKV1TEI8kmaAoO4W6a8C2d0tAB
qUSSjC3S8Vjf82JEJbrDJzq+LFr3a3P46gB2sGeSRB9AWlLIGeUUFtiAZgnKg9c5bVxDoIIdK6gA
n8hLUD5A0+SEg+I0K4H28qU0T2Seb5srw+Jz6JJmEwpAknnKIqulldc/aPBIaPlt4d3DoizKr6hj
WNPaKLcF65a1EUsHrLUpVYtpPj2Hfy2m1sVotSVZR5o1bhrBreRtuCqok/PCNIr+PnBpai6rVlmA
2fxrkfOHV8u8Mh7QWebnzNepoR9VTMNYxHTjF4D2F5C8qAw10cDm2jya9nyoXD3yjdRU1gUGeUlk
v5GKdrbkRlLYNnu/a54A04LeCMdODBGsJRe7Es4GERbXEI/hzqydHy66zjdjmDDLjbxKqynEeQX4
5pYoieX1891bJxSnAEEwEWao6l5n/glVY7T+Oe6IhaXUTLCSIKMQfLL56FQdGqoU4PoGwTnyfccf
8jI3nRnXvlOPHcnsEbhS0cT8CtccAlavDaycogAkpDLLPYU+E2IMdK1v/rSzYz96kyQlWD1XyqVs
9hr3CXK+lvhl9v4PLsQ0Ks+3BGHo4rXYDxkcIIEqUejbOM3ML3mAfRM6TR8Ca16WbyLz0pPAVByH
sz5TRL3oeR3RyjwG1YjNyfa6nZcg2p3aGLZ1zLr45/JF8NRcrP8wgsBBLBJI9aLbMH6h+w58abfV
6D7LzMypp0Eq/L89A7fyDHWVH1/kb1oFOtYYIWF7FtczMrehDWt4qnZOpV5f3h1CJCQjrWrP3IIa
L6VjuKeoYUdoZbRnb9ezPanUPJe8iSj34c2sywy2v+khRdkoLAHy87DUQbW8G4em1aTve0PMA2gI
nVQofc/bUHF03K2a97C3q/5Of6GvhdMB5p2pKIfF0RpVfeZCelCbu7sZeC++UevJkKEXCKPUOWoF
xawvDLLYXNWJBZkOfUmI1LEN0+tHsSn1jzBmeTCLo3y2tVvO14kTVa/0U6yQ1SdZdPvqQO/uOP76
qDuNUzTC6pHFz/Q4H/0rh2sgN+sN7k1fES/ARctDNKXe/8HcAH9i+nUDDzqAG2fjSQgCUvPqOvzh
WoxjhjdR0gzAvgHZ4lk28Ofc7rCmlbWzy2YFgxM2kkjHfsySsrrRLcsNWcPzheTuiLth88qgjx6m
HIIy7IdTlfN0/I5+WyoIqGaDhQ29jCuWf6FqShzsSSBLEWqfFAgwd1Qag2gSbMcx3rZrCAa58yCJ
wIHAvEQ283gK+inYo+zpZSTmS8FHGu6AeMUDi8D4k0r9SLwugGh1F26UMq7+iLl0NDf1eGCHN/ZW
bKThkqRL4ZXy9jv30N4NfdyPb6C/uny3ZMn6aa2KNndHgfZfqMGhfd2tb3C/X6hRMklKx9L8X/l9
anL9yV+hxhUVjZdm4Jpe0FphhX35cdZioAfgRoQrBB5LGINqflvPLfcU90KJomzS2YY8KROSsP/j
IfphGO5AvH7m2jos1WgQISwMUG//wkb8HzDBaVXqUVLvTKZ3/SiwIz9/L2iOGO/zSiEmUzsBZlyg
FhQpSzupqhqjdsIO402EbBLSKAhtgekIrhZFJeOLB5BalIJBZJGp+aws9IpVkczXkDl/7jsNks4Y
10mhaHxtLMowjUJlQ5Hyy6fFGRZ601DP6a9FavQqGR8qPkbn78BH3u06XIjpGxQ+mSESYYnFiBLx
9exkfS8UQpzjU6GtJia2Fy5Dbt8fA3nnthOojNMxoEmwOpHIgEsh29H4lWLCSSvEUvpcn+W2wZ+3
kyYzTwHNkMe7cBv9SIkSndcbVQ1c7HjUnEjX2nNd/arIsSKYz3+Rpesv8aRmRrc/UnDxgoR4xsEE
AbGLWo0Vt8hpKf7t3vx421JR8ki4MBDz2CaU0DyM2AS1Zw1fTbTgrU7blzwVR4P6oTHrh4UQDBSI
NdV8nR+yswfGxhQ/Xiaec9MnRhs79KK0cHOPd4C8BQsrEy2Pog6+eokDnNIhdYnXfsUyJPhha4MZ
esfhVg4aAT1XV9c532+hUcx/fZX+FsMnilzGP8sfU/A4BbaKecoTwBxmhPJJvky6d9SgI8RiM7jO
ZeuluSRnPSAlRkohHQiwjEc92aK1t6YtS7+y7FMVnbV93cXga7N6m8Z1Cz74yL+x/06mXq5j5zpw
OLnSgWVUfoxb196sV2f03Dg+BsVs8VvD7I/ZzAxEArR/ul5vrve9z4Thc9b8VtbsQEZimoxTwcH7
FCbki4Q7SokJ0WaGnAMTYCrOUt0BqBjd1CxHemVLQ7o/jn6swvs8Fkv0is/fGyYU2Kc5pS2SAssT
Jgly6eIQiWaOD193jL11Mtt5VSWQxbHp40nLr1TBzPmuuioAXdheUX19IBccle1uXG0T6F84R8+s
wsIF4/tGwtGhXihvuF1gyzqF9CsdRI12rBs/YfNXMMb0AUfYw2aAXt90KrW6kbvhKDli1EDxsnMf
3IIP592Kpk9hGmD9x4c6VVcxOAGPN+JCiWWE/cIjRGgw0j4egVnStPQwwGI5rEWnW+tC5zyCjE2q
v43EzMfrBcPZQv2ug2AxMvX8bZeyHp3ucsbG8V6+bg8mM7VfQndS/6SODWQtHxUZvGJTAOfZDcQ0
24LotJZ4Z2c0ANlaWsX5ZEuDowUgxTxnH67XfkkWtWJYqMPj1nK/9NbvamdzzCSPpfA+Ltrf8Gmk
VdxAVfKyUB0Z4YpowCMyQ0jP7cVnS4KsLNaSPeozLwzvEV4ocjCUY8UC5KvL1KlbB/IgaNG4hb9D
5XT9nrDTePDVhNnwZr+l80raspZgmlMsdcHhPI5bDc3O5BB9jmnXCrxB4cvI7Gz78eG+tYANrHJG
61xZ0+9y52e7mN9MIkf9co4ETAEb3Z3arPsGtx7I45U5+JGJitDad7scXIbhdigsG4N8T0TZLrsJ
E75oUnKQVu//r2dxUT93grr6/ftdvCc1LopMPqMr6bPBcjCUQi1gBb2pZBbm4amKtXk2d6KKS7e7
EGOx9HCW0Z0EN/OGoZ1HxbSftjUV+pPsINEQgtoILXG63U8WOjExRItGA780miyrLppa+890xX8O
I029H6RMT4onaUZocaj/GeyBhNTxhB5wrsnBZ8FjuCrsnkxc9nS9+BteLks49EJsSUJnU88gclNk
sEbmV8ROpoeIb7pDNNYFcyu82ztyZ/Szp7ikVoyYyM7F7A9gEoz8TAaZ/x0As7kvF18Ml+uRgwpV
SZtjhc3T9kR+Az7RpYn3tAZXSwRmuHJrHCthGgie0jD1T1MQKrFV89D4IsgT5mzzNbgzcjmTNINT
qipMNanVWqF3x50Ev+CrhQIrusoKkNS0QrbfXUceA/ddclPD/NR3jIiqIu9xO25x9HF4izHWYaLQ
j3U/IuDf3vCLL5w9pQse6Ps1P7z6rTvxg99yAv1IofaREsO1Htl6aCFSd7EN3qaDIyIlxSR1SxI7
Oz1ZzbD3Dtx6QCkwND12kh3OFftb8aNAQXLyFxu7Merkexc54g9iCXFzAGAuzR9HNXkdJePnxP5c
27hLcYfuSDg57z62hm3XYLJmpgpG/udBN6gfI7EuwJs8l2mtVwEfr16/M7YGboVDoyFp8iJat4IO
Q1ffN8KPpqZQU8GTK16umLECd8nLTFnI9vLbdjkU5EpttVGWq2NGFJevO83kasShZ9C7OnmcYXWO
B20Nw0clB2SsCLYGchgzyTvDD+DB5eUb9PKBqcyIXz7uUGYEQuYH1iQinBLB3YFfV7Cen213mgtO
UvWkteC3FJGCypB2JS2aQ9VIN8pJoOYX0kWFBrdxLK1RLVkV9G9JVeUsrp0tGKMNGneqceB+CREL
8nV9Hn0j/r+qWUcDDtecCaSgyJ4NWA32WXYPPrqSb07lq+6yF/LYbgqarhae1lVrY1mCCEgPWstS
sB33qtDJZMceDMFEU+5UNes3Zec5pK1s1mBqHVjM/8JFxa+n+a/Qr5xI2iimqVBGGBfwfiFz4Pf8
IoW5eWn15lFu8oOu1itN6Sfq1bj3eEkHPAtFF245j3Gl8VSCtKiU/e9wIrEQDoEzDkOvC1I207fm
1EOjgtutxEPrM1vFoYQpXavvp+pNsV+SAZQQNnRCEZwxXlpQyN6DwiysjpTg1qbEHnCfER9tSg5j
UfSNJ4je8CDZ3HmKlEWa4qk6ehzxxOXJhe9V5WjITjmMO24DX1xxNVi1GsNpez64PQLvmx4ybBup
8fYXHTAK8vacNwYHvQDFtlQYW+6WD+1LdUoGYTfIRn5wE5ZtvopRHk0VgMTvFJf2zzmfx98REDQh
Wjkx5r+RsftBXt8Stp/LHmpY6o+udUQ52IzrXnoTO9pEV8EGO2HYux27HCWoEGyHVV8ad8IUbI6E
z+LQu70kZFmHqi2RSrM3N8UPFxobpfBvv9xWsfSJ/wrV9LEDLAdQzOjJsu5JuOtEW9RDCAhoXq6Q
pgpAymPWf1rYr7IThmOP/yVm+jWxKohi/T99zr/L1s3KQJAtOH6a9wCHl+YvF1h0TLq7nWoMZ2zP
OAdkRzB9o3ONqj/OZrd3adqos0r2I0Z0JJ2sNz8encvgA2BZQBnHUybJlyuMDepKYbp/z8uYKnAN
+Z1DUDddExFDmC1X2srP1qFTGT11YgIGAL+ATqMhB6GClYKkIqa2kXGNcezeKIxeBn9Xb7HiOxVN
I/SFrDi4aAAslXDaqYH4Qt6Cb38JAQdZk0KUAvMCEfHd+2Qpp6UEQx1NLG1xtiv72LFLj4AenJxk
8JQ5rtLkxzjhGYIsUSF9WQmRuoJsUkK2tytJgNROoGdjuBgouyZXpglSA2voH1qiUAsFf10QPWdE
fv7D1fuIsLnuUaaUDEGCw/idrJaYPU/2w9O6ELj1TZ67GMHwk82Ekd7hdIGMHY3TWkSAP2GxuT56
bUwSxW9fBgiDDZlGok4aPZCf2kUbS8lwmQX+lBqJN5Zn6hKZ/uuNi18135WN6JLAhHtyd0exfUXf
dffVs9OazSthUkFaYU12Ps0K9jrU1lAgkj3fGFbVe/6aB4md/cBjXNqrDDP4z5pWNnYrqzHsawT9
lz2Pv3pkXjwwvqNBNwZi1Dv4eYALDpX5Z3jNVZblTEYH7stCF0TPOff0giSk3wuaE5vzMDtaXKyu
DcrCh9NsytZk6Q4DEoYTrDUM1X/oRTaaf3KmTuHRhBopPCR1ISGjG1uOxTmZ+4kmqOygMi2wF4Nz
71ASoHJihs0zaXWPHqrC11XAehrsAwifdX5K8KetMtXqGv2z2Ty1O2bxkCL6Y3JG0yg7+CXj+i64
Ldp9rJNt8gW8ziSWiLBma8OXXZMbTs/1rEhqNLrPlSEB4tqWXazlWk34zuvj9QZfy1wLfqRPxgFV
8VoZ5ergz89UwYx2/JYU/HDKe8/Yl7AHi35QyCn+X3vX4ukTVNE7wy8jMjrM6U5cBUv3DNT/XDDH
dxtT8N560XN0tM3ea4oZ7FXMQnZhD8xpQ6wveZFuVMrEQHPL+AFhT4EgRzUdrqUIVi0/4XkY50Fe
z1YWaMHDmJ5En4jv/R4kc5LbqtNmsJUGmRlLjAqXZEiXiPInCN/G+qpx9ZrjIAEDsdDLC0KmHzTq
KPkYvMN/zD1h9NMDF/aMTwH8xw90E5zPdaE+hnADYyO2wMDJ/lCtorzyvAwPSGr27KLlACaoRJxr
AH0fCXrmwahyhB+WbrwlxJ1tK5TPAX3V0VmCh3r2kQ4Mttt2l9PhS/ODcVrqiT15uoYnNEyKzVIY
VrFBVIhUQpMRZfdh3eTQEAtomUjo9+S7i64o7MVhRJKmS9IGNGeEK6jbF+cH05XgJcC2g5cD3jj/
dl+dKJHHcCLQiPaeIi/AIaIhYjD8IOAPLpsDKtpob4c8SW87luT6FXIr8A0F4N5HlXN73OYNbZuJ
t1IMv8kzdojG7dIch9lMiqqPviNlSO3kSq2fAw1wwKJ6WlK/F7vFIWgvZgCKUkcX1vXlPRJg9K8O
gmMQ6+XngqfjRNsKEZLLtHdICpfNu0hvGWhT5yKIU/wFZdPq5DPMsjIUnRh1XE4k5v3WNa2vYv1h
qTiSZNrXg/BXHtZX5qxtF3SAAkeaAKr5rHzaZKODcgdEqg37NG2COfq3TWByBM7UiM26ENMzThHP
QyfS6sudykVd+nG2TNYE5CnB+r4j2uZ1KBjewNaKZymoWqJK0xZapzGJRYFqJdH2Pu6IkbUtkLtJ
1yoxHqgsPDgowhDf37nDTA3zEF4XhkXTDWGKs9nPID/j0q8ETJ9AJ1Xm3GidW/Qd0G1x2Rc+qF3K
e6DMWystPYYAFzpuQ4R3EvdoKp7lLHtrZ+QPvOsf6gk7i1+CYVcbra9evV9x0MBMK092cQhoDLqo
+Avq13aoozQo3Rp/3kHpmQUIFfZmyjrNOVryiZO6liyvcoxTcvvaYr3ysW7wVwYMG3B/POADJqWd
zJKvWWpLtq14woqjpVMI/NCg7mENhlGfn0QxbQqbLw62o92yiq9wjtbKKmBizM2+Fa+tYD912Mhy
Z5WbN1yD2LO84XZS33HueXuxUZJcwA951zVp5NNxcKv1x672G1J8028YI4s79XNjA20F+p/0lxjv
BkN3ezXGM/YO9GEtlroq/a5p+FxzzVwAtlGz6iYVKBDwQzE8ewuB4VKrfxk4Uuo8GkuSgrpCsbba
tLo+tl8bxn4cJlocolSjBd7LADMNqu8BMnBQKIyEazJvFr54T5zWCLCDxAbMHs78+Tr4A0moXvxm
Q0Vo48I5G8kEZwul7Ai3NTkdtjPJFjxWmtIUkU44c2MhsanrzrOIMMTmLBFBpkdgX9TjSUZevOL8
oHw/PvAiXQfiHeNW97xBiORNFUf66Qs91px6/s16Y/pwrLdKHwNHHWEMWUBBXE4q7GdxcvJjcJiP
eh/RQzIKHD98wgfuS3wgoy/hBsQGu1NszB/fUhIUS8wNPLT3ux9MynxEEspBpAYHmANw1unbYHj4
5DnDUQ+7La1i562U0eXv/221DgIfOnfvImk4cmAS08/v4WCm9OYcr1gUHl8O6GJNbrkjBYKm53mh
9GVi8WygRxQG/27MW8yvVTDGV4fIWxph1niwj8NuT5rbXkRES93+Q8LIqhmrCybRPh9dbKZJlcH+
KMnc3npudHZAM3DKSmo5wyildAy4wiFMlS9GPpUZn/bw/6Tfotlvf1RV8HtSglJOvzr+SZxGQiJV
m8xsC/5y35toQ5+nnZ7ol2VJzQQNBYewlVnyVh66pzAk73HfSkr/Ty0nHFg3qE/5kKWBTHeTboAi
sFkJaPaxRJ3kVK9j2pjwiwAJo88tL0TOwuUc7N9YBXtuf09rDaU8XQ868X3nZBlbnCEbx2P3TcmP
xhbvFoNe193jzVv/X3GgkXQb/jhhUcGLGP55oz58MSN0H601lMZHQdR9O3fR/50GfT1JSqpbzRNO
+IzTUnRLkgTkHY2h1cZvoRpQe/xps2hbL7GvnbQ0ErhAboykosKbJz50jjwrNQnEeMeEB3qbKyYs
EQdiChnT554Nb9hRVHkOYOFuGsw81csxZgnvfnrFUgm2HdBFYroRoiA28HMnjwRib8bNhqXtLN/2
gr7reR09czk3JeuyX+EDB0ivQpklJCYcN0KJecOwrwTjpFwYYvJIVwOh6C3kWsOLl4bk978hbi4b
5Gq9VJ6tIxHvXZTdNF7kWpqucL8KavOdmJPMg4fPc4khznIFmzlxJXa0vsSEVYPBhKufxTRwr+5n
+2qGctYDsG2XAAtw2hkkMNYZeZPp8eBTtT+dd4kc8DcHYCvVVaBV16bzChRzty6crkQijmM+YXWB
GuXdPhmsX1eMobpJTZw998LlYMY0HVH6jKZ6GFTg8xoZR6MhdwdDsQSfsBTRk11i3KtbZIhcOYM0
tbBO4CtqXzSjGwvSgY6JfBTTDb9dmjRLWnRA/gfsAb9SWs9H0Ua2xeVelmgykBg+ikzvP6rmjqvp
2LLCYn7sWDRPiz3deob/mFYKvYyk0oyTwm92/9LKBb97gXjswCynFtsEhW8zhmgqgYc+9hMl/gxW
DCZIRPL71ALKOvspReTdZaxFkWZw+C1Z+97ahlZH/CEKPg2uULJoqJLRRwfpslnmHXsE9q8vEh+l
QIqo5PdUThkKNnfNN/UDZwsTBeJUi5e+5hABUkfsNxLoWdSLhgpgWEo6zuPb+rj2zyZZf/E9lurV
+/PQsBtyo/bMP9PI5qAQnxL0jwAnzWRO7GRySIPnQnz/rVGdkITU+ZHn3LgMEftuVhhekZcUKdJk
MZIkcgAitAwiKg/U8pshs3qDUoOTzEi8rDC8PoeU8ytIwoJ1OU/1xMDLiOQZARIilE+n6jJJdlFD
r3jN07TtOh7BV9T6NV6UboFAtNAGFr8WSbBLoxu1TzxYMa7eWfZmIvKuyZBRFTy8ogUyBttLhrjY
MXfqJEWuT8OWs88Vw7LUqvjfws7SCiEn6dedWbCjahjR+IbIzDTKimy2Q1DzJCmu2vVfpwRLMCn/
52Yo/lMRqOZNO7YIF3pc9R5GwsWvF0l+6nf1cTKVz158Cg8IWT2bDeeOnCEzx3rq/GzYYbKzMOET
jSjndrJxnz0Zgmo2Q5XfdXjZDdVoLd7XnpmR6XHAPVpDRM1kj/AuqADaBNMal6jS0yafF83llNhm
JfauIknjR4JQ06pSDDIQaBcq5mje3xoYZeJ8WqSfqPkbJGXs5tCgtk+c8Iv/fW7ufKnaSB+16Q/s
uBeXobSRdVgkle2NvgXPrxDfTDIvgq+N/4lLSMijnl7MDhhyl7mG2kV0eZsfXGleuVe5cblzgPVb
M9hQsi3JNpf/64M08I5tu35yLHWmjE7f+0gDAHKBbc7ngZKQjEEA00xe5krN1aO1sKM55eQsXGB8
REuJ2BlU9NXHqYcMuKGhVRUHJ7/9GVsMeqeKvsinGaCRMEC8n4T5ko001czqMZRACL7/PdIoUUAz
oMV07keEoJTsBQD7BdtHCFAcN3KgiEGzryMzrRgOUSUcpsOvcvKe9oCgilqhpM5oAdRdaW+rgPs9
j7pTMxR0pulMKJ9hhlYkjASWW0rf92cM9QpHJr6QgpMhs06PXKaYOrjBc4UYk4NQqjcC5AceYAdq
NEJ3AaHsn3/bZWpln2rzk0nE6nSYXb32UWxT/TYWrURuACLfDO9Mb/YiZCL9jvfOVAH8Zawip5iW
UClYg6z1o1XvUT5SV7yWT/bFGRDrT2H7AN15yHeRdy01Xan5/Y9aCN6ezs1BhSuK9+yWGh842V6K
TjQ1lVp9vBAen+Gv0LJu4LL4aNr6zV1YbpPWZWJJHSHChR3iBzmf/fJnxn5iMNLDk+a31rLj8PLN
wE3/svDCO5iMCyzmK9yIs7t8ptq+2pElxPpw3eEGJdYfRJ2srOO09DMXI9GLMEutGCeIp1PQV2Bo
iKMB5t2mxtz42dnk0naiSCjLS/KXOr3hz08LAnspZtR4t4ksI6t6bwgOuraoaxi+g8PU7J1rs/Yg
lg+A1mXutj2DsnYuzgrz73CnVnNzuBGfp+zJu2OQyHh3NI5iGdoZoQuacHH5b/UmXoUobbFBglaT
tTorvr7UiCbyNc5B5sTC8s3ROPfhDkHukEumD/0qItmpERb4YxOhCxjOxBqa1kyB0ISZERLmZ5Kz
q5HDl8JJHqWJ7oRhmgu0xm3azVVOpzDc6S7u/ISW6FHEJE8b/Y0f5Z7pqNj0rvxJQX22ixtfAV1u
pPGflW7BlZjuy3vW3sV3z1t7IEC7OpjT3+hunWFJCcJTry9Ctd4UPyCh4qgSlexs17+0Lyjqtw3L
HCi/9HGKgYuHWt9TCeDOagytaKWL7H2yinvRgve+wKSTIMX900mleuoR0p8DMx+yfXLrvFaT7mmm
IwhQ3Yq1P3BWYHKnIHpEavj3itoAJEwujaKOgaAnCLNrVI+413p4e/u6QvGrGW3ZsgSVFc27gjQ8
iQ4oGspfRVMYFOuzrrOuRYuDyGWkzpY3K0xs5fok2dvj2XK1JPUmQAopsMtnLm+F5njt6k197rWa
Ov+124GvuRx2FXdFxOlZoXuYn9d7j8N5w94WYFFR4VYiDK/2BvjWV4fHt4e4BOme7+bSJAUNHeJT
Xzo2v0Rrr7ltMK2kgLT7i5OsBeSNWqz0r6QZahsxwykqj7mobrzjDsPo4Eel8vvDdOSHygDmlhGP
0IH40pnX+xBAx9GUic1j1sEbwUZob7jbrIPd6EDirsc6Paism9IlbD0RJgtb329+WYDLg9+dm97A
DSiVmN/H5whaehAMQOvGNc9sIbjRQTwnRskcpZk+oRIGnkf8qlqRY3g43RKNUtHjlpJhXMnBhGFh
m5q0Y8wzk9oNpFsGegZ2Y6E55QaId+WLPAMmSJZDjgCSmwlkuaFqlVVJVtp8VmirPTSc7WW5G92S
PV3fqmmon1YtF4E7ef7ZVWlyY0brTm/3H5TXT1wNEk+5Dfi2eZ+3uA5D0VtKZklxTLh8b3USgOvE
kct1DyuaEdpWOpi3+UMGA8WPK+lh/TfJPprgTSIdbFMHYC2Y24QdAllGy4tgjlJ0cWDQv2ScT1Hz
HusqJXDlJ+SoMtQqrv8M/f0qnYVZmbYRj+MHj1+m9zlzDzQNukwCaw23ecOx8O/RPxwl97JWD5vm
pEH6gv06o0tNziCog+F1nfkhrpIth0nlRbzkFGr+jg4o90tpNftX7ANYVdLHfJ9Wpc709bliRzX6
8R2+WOO3mVyqOBo7vBUhDQqnIQ/RqNfPrFRh078huK0GV3Kzkkyshzl/6IkN3RMGo9qZRWH0TFVA
/pq4KLKnGWmD/k55IG4Wdy9nzLboOxmzsH36ldczjyBnzk7iGmkZAjzr5QshCBjypv0nfbyfGd5w
UjR4VhbwCY0v+ank7xPTzwfTjxmTJxDaAW4Q2wI2s3Y1cagWbXAgyA9ClIKoj8RLTukRmTdMyt2U
aWB0ta8iBTmHBbHwH+w2QWf443t1DevKt/+cALkaHGbZ0D49q+77mW9+QBtm1lazra6L6aobYjPq
swam8OR+yaUOFXmynqEuMQoevjs6RYm/SO6bEM/AvMAsORM0wocdvHOSvbYyBzSot794Y7oum9dO
0Lm5sqRUS5fFCfNjt4gmmwzbP/6DCiZDzbnOpGp4XoSluJIvxM5RHftAoxJelfLFNDtxVJhphku5
lKHktYQmAfzeOCN8xPwwa7P9zj6mbDxwVcU+FaE8eWsDis1xESYSzBSAmvMiWNdlJbUCZdar7PqZ
s48GIhngbbf3al6IZYMVJ+4+mq/uP5uSbQM6zEM0Ba2CEuHfchsi6Y+PmWXVDC+SocHc13uqPwaw
MGDz9W1aJ7qHxXISJ70PuCF+Z2e/r+KsrNP0aZXQgwuqL8HCWCLjWbqQtxbdRdZYoTCnVA6xQT4t
KFIwAD2/0yhV1HuJF3WzkCsjoY4T1iE8vmHlNdB34YPiCcOah1AMT+KdGVOPlLzQPbH+pRffY37z
XTWfSB8WVz4fdsm/fw493iu7Mn8troQ4fIfNuFEVQaGnI8YCu7mvm4XaUJS6KlNiSxBjagvouiFY
maDp685N0yFFJI/2p6apSgEX5i+cO0ZaMaZ7KuLhIk8eBZmQt5rFciz71UTUEZn5ubCgYwIrvG4M
kIa31eLa3HBjs6Ss1aOwWrxCW96tzN+ciTyExq1iSbNmqpVhACmVX9qG615BmEeDS3lsl0vNUvfq
jHuMXXxXPPUDCWhX1nPvmIMrdsaa6zQrm/ZKAKiqENK0azwARUdsjdntdvVft/Or8CSp66ubPrhe
6qZFRnhaisZOOqyVnozXS+9j+KVWaz8lLl2xynhncfuHGvvlKFE9w4egzXRkyTmDSNPBOYOTTWrI
oL+XPkM1VC68vNY+wnO9w9rE/NI1yTMa7af3sIyviAJSMuUMzN5EpfdTegXRoE2sf+4fVXMT+p1y
0oVo1KOMD/98A8qJ1c7rAl0q27xxpELeV7BXpghVh9WCkebnvDGQ+4SCKg44cPXN5zvAj/jGSnAL
eIQj/Jc6SKf3CeVhiSPmQtbL029nIF8ptKFA5kU/Abln8ylyzhOa8Qj2cxZNbRZ2gWBx088I6vJ9
zGTHGWNVr3tz2Q5BPqVRvCsTh+V4w1DnLQ1xyqiDoznmU0R+VoiK3mG+xwkTF05L1MEGX6cjfiAM
aDx9+1Qw4n1EWpVo9Q+T6I4neNPJQlgFWzPuLNDHElP/rpSw9Uj2Lu91d6vOYn5V6ICnJfGGK/1P
B98jxSGiLUd04B0XvM/Br4/Gby3CmdWI/sa93niSWg5dzT3ktUovj/ieoZrgpKQDVnmq4IvRLDOy
5w3S4hxAeIyEWBumLsepSxHCn6y1wU7yLlEpMOcMoXgtuGtkQ2uwMPDnDDzI4HiyYC0LVtyH6pV7
kHeAbGv27jlFIrbzAkitWdsIpvHirvhho4XMAuQ88jkcZrmK5tW2M1VporU4KOkyQ5ROm8OoLrAr
kFsDaxYSYFvwElLJcKjq7FlbqmoRPheKY9uvhwJ/ZtrccKc7Yo0MFckb2mEwMyRiQOy+bpCY82vq
MWgb6yINGdrR6jqkg6m9rc1/FBbCBx1tdxoHPDDHH0rzD6V+Ap8vz9PT7whrSzqiRMzCsJ0yAjCq
/0l4c1jd5A/YhavuPEhE2ylWiMAuKS4dX7jtik6xGBlc+m2zjqk1jZzMB9E1rGE2JBZn8gTisV+L
+PBNcLvDJw2AU6C52NJ7X7YlpefwxmUW6XQDrPxcydo0UCnFe1o9Z6aS+K0fme+XOhF5ykv528r2
ynYaZfF8cpVaxLoocSgErrmi0FRVB6+YUsPxvTaf6zq+0PEODkRAL5wpIY5ZpL4u8isvNv3Wz7Sp
kC+ja75ctoVqjnZUMdpAL2LvL+TtSp+to+Ot0zfjYRYiQBlr4cQyUxXtdzox7+9VEjBVoHf4bMnc
QxOWVl5vlD58i8GZX/gb0mE+jgzKS+m96ery7SO6YXrKOwuGV4MGicX3K9EYtQZLbwazDfzyUQ4A
IhGpt6k0kY66qwYkdtpUl9SPh9ICvZKJeyqaF/MejDLnu1K56K8PEQk6OyDWsyxBSvxS7QhBmfYB
iCXGHBdZyeu34Nxl7eUDiVJ1BGULkckxzZ+jFiWy6+jBmlaFCWGVt3lAp7+/G7wgUX8ymxI+8VQj
L6npwr+sda/0iZyv+kx5/Oed807U6s264w5qbaU+Xpbb0aRxLUF0uI1PH9wCBjg8K2X8+vQDZd4V
Z5kl2aKI6Efp55F9VVq8E34KpPoj3gfOt0dJkIRq8sCIicY9ZbG1726u+i70F+rkkyDdkKCfspUR
ET2P/RwRPNak/ag+PPRZB81XsqsVjXgjM/PIBP2Ch6zekGdOoAd2wDGF4D5lYZ92QbCRdrxBGYBM
ZBJ3Gq6uN7HuRjOALzHVYAFHfnVv5mMUHLbSTlvXT7+1+ZD+cNeE7BP4XQHZsuDoZRu63VyJO6r6
roQWE7Gs8IzDU2oJ7vLsBHFcFRxKHWjx81Pzjl+8FN8qknQEhWTQAIYvnR5dqmAWl+82u29GoqFn
XMKZLSt2xFDLom9pWNYcJMvXuychvqMD+yzTPlh/eKbx6oEBWdq+MZ/FyXdZE+dVcTs/heaSy0vX
wKTMe+D0/sH3RXhdx7anaH5+LZGjPz4oxP4KEb++b5Dr0oYTPACDPeC8yXCy4uWBCplPU7ulC0sF
I/jyFmVvKltzfE6bdcjfOdZC3lmjvELRAeYhG2edGDTCgAVvNZaIx6Pp84A6TbQ1fkxyGqzflpuT
2LO9ghRmkopuaC0RofgYEL036RAI8EiohoVtAxf4Oov1XkNvvG9qLNtS8aqelm4cpbg9fEuPQByU
bA2kN43UpbL9V3CY8JSRJtAa4DULlxvQWhR2QypC3KFenmskpOG9sBvuzDnUwiY360boXi3euHMN
bCMsBeS5x7Y/EsuWpSB0+ot2qsHL1/RvGE2oFraBOWaL3AzYoWG1+zuOeBCc402C4IXrleAlsiXK
mdPwmym5/cfB7cHWpz32Hq8dOmp6+Nxo3w+15RgSxFWC7nzVj1o5HDoentSilkGU/k1l7lV95YLK
WPlHZJFetRO99KvDmcT6e03UMO1MjF/Q31d1azUES3Y7jebI+xWcY2D0LRkWeKBWz4zgC3vRz1w6
kfsxZtvSX4DzoSacKyjnEw7hSunnjg/OL+mw9MIvLxCe6V8ZC1Z7e//XIjCzUivRA8pU51jdMm5m
aGCQJtyrCtWC+DnWsQ6DJhLR4LOIpkirLNlmGnTW0iodw1UXBYy0hGT/0CpW/TMs2vWgLoe7QhA+
QMZynDB2EdgDBJqgWmsGo/r+9oC+OWDoBc73uEeZgNNwkp+c2sMbl9Mbbwrtj8zxRcNwvnOy53lu
9jMMTxY5zeT1ZO0erKSu7bSNWIk9rByvR1EjqgF9Rs5/GDBO9w2CMGgakh9KRrW+jcT/saHviGH7
JFE8Q5holi19Cjs0aSg0EO2nNg8Rex+UIK19N8+Q3vSPpjytdu+uj+Wj/TfMy8+Gl34ti+xzUoYE
ao/dBZdlzGmHXuP2vVkU6xkFw2PCqzGfokS1sBs4rZ16kIhhQ7pIYL0hgA1RmhiA3RY6ETHv4wQm
czOZlJDISNjv/NX7MouzpnN5CPCoKpk+URRrU4kA0yXrqikBVwZezwHnEX12PNjOpcvOW1tGpOTX
jgA7b1U0cmswBF4yhcGwggGUsickHQNT3VKUuAjN9WATCPzIL42LTJCBj09hTKv7tfqdzf4Ou3sb
lEi7khjQjek4t1DUtRvykrCgkLJksEepIpGRjBVwQQKmNDYNk5YPl69QitRczjuCn07UjJLiehlC
Ri1t57Woxs1PiBYhd9x/U8gXaVM5KMIOsLDw4NRS8NLYD4ji1ffvNeujxXZ7S7VR2XBZSzjzUkpn
bhq/uWHUyM7pEaszMLDMHsyWpLJOXAAhmkYJh+n1pOiRc8c+pJIEfw0tzYol6pXaKnvC6w3JY/RH
QPqc33Spj+qwesejd1Lat3BCZcGUPTJpvmIDOzCGhnNf2jFNAVXYDdJdYGEYChhTztB5KpqBBdUd
PCmMknRifqU/GUd4oZdD2nlOj/dtPdbmd6QBBowgVF+enXErjq5T3jiirICKfPA7bilarXWi/7kq
OovY11Y/DwO2jR5tbJe13TJKmkdIDtKke5OXeNSemMa7LX46HmRC0ebC01ninv+fMtl7++i9ODhp
0oI3CxdpH0VJDpG2HVsWMeECG1gwr/5e+v6xPDMIEiEqlG6D8GdZvF40ruF96jJcNu8B9hCbfvvQ
4fhXpP9DpNvoNqdS2WLeinEBJBfEvKyDrt+74ARzKGRm1I3Ybv2vAPvYiaVSmdWNyXMGOIVJrwTn
X25bVLPW4qEycxo896OJLZRLP4S2R3aA51tpZxgU3upO8uFdCzayzl+dNOE9ttl2Sdmr75+LN7VE
52s+3AQ1mp46zqQPcrZF7b3IXQdpU93tCQDYKaARKdKhWlarCDD/jyUlH9LKRvink/dvMW4X93Sv
Pw2zRAXbDkuQnbDgBRf6Q+PLXTvl+PA41UtL4Gs3V03y57bLnMbjO3QACA1gQZk1ws49WxNKq+Rv
NuGxP3Lrt0r5A/MijxvT+g+x88cI8ZKx7dO1gjyi3iMt0RQVQs8gvslagAhO3CKWRpzaUWQaq8Aw
E5gDihIA4IceWW/7yqluGG+7TwtB1co/gYJbYeqyVVOnLn7Tb3754HU0hAUQXRbLqHmY5Mx/+VEp
/TT4q05fIcsHuZOz8Mbwkx1l1fueOuV+paZVObZJbony4L+AvKOxojWjuW3MfZZ7Im01bgvAliIh
pkSJKcNxtwAykLCQDKrBHyBs1LlZq1OwHHz8X6XHOsABaCG9Sa7AKP/xcLExvd4kv4iLEvA6LLrX
lMnGLQsK7sLprwclgvgnupPjHf4NtA66j9lq8opMNqqJHoALIRNydPGZ7+X7GYfFSDXxa06cqiY/
pekQfoGbplHZO0lPsMOERH9a9tkQCpFtBzyzpp9hBboNpjQfsLlUy/VZJszI0zqRfCpufgBTPRPv
cni47KHwpDS3qy+mdoVQwwBdkinbKux85HDPu8sU4VF1U9i/uC738x5MGpyuUPU5AcndLhXvgW19
dZNRM67NYaSCKnQx8PJ6Mkv681le6R0pSZn1Lfn4SrUMh2yQfxQPvTmr6mHanWMoOGIZIG6JdWdz
iBrDgODdGMG3uy7X5v2AwqIDbe+reFBY3o5Dez6GlMuJhNk5+chEbAA75hewclpXxD5eZ6SA9X5t
e1bclxkM01CAAiugWMiEYW0gQcuIOyFmD1q6V+qtS9KitHkWTHdzZk4rDD9t6sMimiOftrEFW4S/
zaM0RBpUsCs1hjyEfh8m0Qf5UfGq09uK8r7SyNIIlkQGAut61x6X4Lj78/iHuMaZEZcDpQWm1/MZ
Z/o2vZBi0TJ9+zeAR9tVd38HAhVxR1Q5XpCehu05rEoO5Ss6OFJFU8o3ztB0i3ISivBL35zKQu96
L8aNdpTQ0cSZJOEfQDY5I/V6ChhAf1kIGCC0ffZwjwD+tuLr2Qfch7CbFrPTwRdVjh2489Y3sR5Z
uXxKyXRxvUr64HhwUTkEvhehkZ0fyLKIBAWy8OaUfT856rI16Uk/AOvSRp89HemN6TFSX1XQdhTT
ET3GCJEyCzkNGn5JyPPCLx1hdIVRcWIEhdZA5e4/WummojN4JNNO4EpMzOymdddPNs9ZHtkg870u
ImWVxRZCDsZX87j+lQU4mZgGSlHH8mxjZSwcOS0KaTwPOyF0OOVwwONpGaq+Lcv3X8SLs45KNuWV
lAb9toRNpOShWEFz42OEugWw1S699WPkD5orkgniwqMULAvVvBozQQbgInwJ093sRRAheJYX5bYi
WGZm4eWjVyy+3exnS5S37Kkqz2Wo5QGy022Op0i+DlCocIEzmUPScng4PBQ42hXCKJ4wTCJqtdtI
FN9yp8KlwAQgQB0r5v2Fzs0rB2uqwrPmIPD69lhJF5zIVsV52c6nuQ2bJzicx0zFg2GnfEE4uGBB
pYNyWxqSZhZjog3faHg8zW1bVmbE9KM/mMrvERSnEHIR5A9+zj2BV4NTwx3A/oOiRK9WtK0D4Xy9
ytfi+eNqD9GOG/05BSa0Yqlnhx8ziL6+89S3mGoPExGtdu+gIVuPeIWQ6QvYTA22ywJ4r6SvX4v9
h6KOqiow+wDGIq22dLPA40ySJ1ZcC6vi7ZIVBZMHbYaJAF/VUCk8a1mnaftgIEhNW9831+8UhL4F
ofvtcmfp0PCDZRGA2jAEst0jCR3qmYnxJlRUS043N1CfhNTMhgqDGYKecz8vSaDLv5PKhAeYiQuV
jZ9YHMSSVapYk7NoHhwufFwtPEPkgINn3+eoZy79mzYzIo0TO5K5e36c1fHlkzJ1AmZlaQQgy5j8
xkSt4r4PKdfuuE86tb5X+v5AiqafQQNQVBM6gmtKtTEn+PJIBYXmdBlrqX3JaY4aZxNlSFk+gR2i
qiGjN/gDaYDrUpNb4FHnhxqK44lM88/VI2djOAGgG9IjUO9+0Ap57H83h2zSINs3g+4vUg1KUrlZ
qjqjyRZaCiISZ3WS/FWWU0Hfwv7FxhLjvdlSiyk8UpvrzA5l10GprGisJX599jN8JvnK9cg3A3Fp
g1ONrGHzeGWfQWFdB8mi4dtI8mCIM9I6OQEOhAWJdyHUHU53Ir/qekYczbYh9v0NqIoR+U8lDG+s
N6ZKwFyT5rkKI5CXM8PiC3nyvIKNIhsQ4v0oLTIWmN27Dah64YShf/Py92pw+JuCY5ieyOm6an6M
jYvbD5SC5etzYjv4gUqm+EdTX5IyNVA5l76A7QjxfCM4Vpdmv9h6e1YzUyIL0FeatXpIQUskPzFR
fKBXBDxJAdlvDPy1ol7+ms94IUO6hkWLVS7uuIZt2Q5mmO7gNeylFZIhZlvasY5zDNNAvnluHQ78
WnnBiV8L5SJ1XsshivKLcwGr3tE8C2W6JuXCCi4Q7l7Vg/vE3cbSpfCqnLYLzl3sxZnI/7GGu/Mh
n5NC+zlyk/LFSO4OdFJL9CkhkrQH+OU3UtZJYpSVY4G/d8oJ4RolJ5oDOr2r1DQeorGx9gHiDEIL
2oTeW+fJz4jfR64wc3njRFQf+dxQgQ3EiGzmuCsJACKczJh+ntO6cSswruwKBH5WLvMWl++8JLq6
DGEoL7WWz/fzPhkOb77AM42Ey9PUd/eh0cDiRZ/j9LKyrw1CDI09gCiHh9Lv+659rYi2mbe4OiwH
Dbi3TpuTyw3Ntgz/Pj0FCFEPnm0/ncjmfe6vXF4Y/SdbLVIuEI7/yw7I/PwCpkWJO1QfmWXh3hYm
lSHf4a6Z308HDmH693oFYwRnRi88U34LmBH7NtzpE6UtNJd4NcmJMAvTgZEE6XuuU/IbnjLQPPLh
lruQHQfs4g/+k7K61awJOhgD3n9oNkYZUWWICUzKkHTR9rXDkDP+j+h4WfaAMcnsQrBthzv3PXee
PlgRHwSss330opcEPVzrcxREeC5/SbIp6HzXcnPcNJDXstk9VqMWnN6db5aA15CZwjY9NfzQryCM
csOGuOJ3g+eQdBiuwHR+by6AJPRQWDQik3YvTJF9PCa9mfOOYd7tBbZ11YLE6wubJglT/a+OYpCP
77YjHzqen9EMxjPWq8ZclT1bOrZ12KuCX1N0VOgN4D70beoaUap/BZFfaukh0FPnLHfit2kutmYm
rGQGQ5anWP0Zv7T11l9pqJSxwVIxIctUImGaLUfT2H5zHFky7strSIZ6SjPgSLNdppiXkWwab2/L
xKsJ/5khqhgHixIsQ4XGT3v/A3L43Sxg9k8EjwDssJsPZ2FnIpL5iqgLrDzs93wsWldE21rYW4Fl
sN8GQNrS6hO5NKNcM2Jt8zBS8WgWraWiOKupDRGcHyUoKJG8Qu1/afXKvOshWC+ejhvM8oddGVXT
su6j/rP9nDfa0fOl5BUbMtjFpTkvmaF7qmW76sPoBz1EGaFD4Tl8bdhXFmv18GWlCWCXUzlSuhml
AqMjCZEoUZUZTAdc4TXKrcXry0ylsjXykH60Zzr6o9+M6u03uTdJ99SVn04iKJq4UxNq6IAWVrnc
zFw2zl+PMWk6afztNrEXCRLLwMQji1pcrkoBmbnthZMgA06UrhW1W3k7RnCLdHRt+O4Uo41u+GB9
0Qs8tXeK0vptQ2Dr1UGncyXRTt5VxXqH4dj9VcNSDEdv7u/QkwavqqkAccJ2UVvS5P44tKYifRTD
4epmeTHlFjF+vBHGw3hDWvEZPJkZNlZvQPA+ruPkDKkY2t8+dp94D/x/iO1PkYUbOK/uaXCYe0t/
AivRu8/+M8siMFp79Q2/fXhkqLlX02eEZJUxZi2aqTPKA2w8VmcrDUXh3PG1LmhHd+EAi+TET57B
pZuCHn+RhT3SLzOOlcSMNjvVLcq2U9yLWN+Vqfcy2Jpq9Z3JutAVGCSH/mC1OsyuQhaafZxq6bPM
AScBZq7mS7MqNDJPKIsFvnXu6qD/sBaE6sUfyiOBD7Z2fmAs2e7FgvAHRT0qk1MQgtXor03LRdKF
oBym+IOiyR6tZH/JVSD/eoBYCs8PmiJG645PMS+ll8L5ecFVt+pV751fhbcaCcZydcDgycFUit/B
k4/3hI0aZ62KwEak7UlPhK9nX2aOUU07gOf9PFNIeX64gipGMs3dpb2ggI6m2DlGPPMHAmXx+y8T
Nz8fHyrkINNdklrkZL0mON9CsPoTMivr9CtWU2TrsMfYpqVMbHRxzxMwWnTC4aRYYmeyAbi5WxI0
/EICXmUhjKQPr9dUStr8bay57MxbzJFyS35kSrsATbxqP8GkX8qG1RYGXafA+8L1taNgnD/al/Yi
dfk3CshKMWoZWNrwupfO8krTISWXkI3FO74BYzpbFFCvtvfhW8KL7rzi1r4zYTqptMv+x2RLP/mB
cHjbp7jeQXi6O36HZizHj8hdhh3aRoVznu8vVy7VBtwrTBBZSnbnZR1bb3CzFr65vcaWFCbNqbSG
qhenQGsJ1k0kA6EIVx8IVM/SEAlVd6GYvFh5ADmI/CVV+VbMJe1mBz76dKKDxfKwio3rARkzlqp1
Sdg/TWoXijZCE9AoUlILP27grE/IIspafYvGBRCUliLyxGzYce2IvAK3Jklt35Uwh6S2oPt/F6OJ
3mFLVPYbjuy4QKkdxdwbinf1gT5Q0D33kJtZ97U+TfNtkt6qm7puOwQmOvy3irF1KA6ZgS3gRwgN
EAgPRrAo0X3ACQljz2jJ8yTx02xTis7PwrJleztMP5ImhLEc9/sVGF3ER6lCi3i7o9y/coCvu4CU
u0yh+L8AMKtHtTNTwVJv7Jf0Ao/a6pWYDePlgh7HYjl/HJ68ceYO2G8sc8XKtN9zn+4fTy+kpaMT
juuJaz5r/YSjnTBJRUWJP6nqIHV+7Zxc8Y3IaPytySZRBiXFRLw/vVtEO2EwbFVwKDFEy8gANJyS
5SBGWjgUU76o9SLPpJi4ecUs4cb7aaGUq6OhlZpjOhtQXI6fA39OHlxaicMaX4gXC6kAsAp1k20j
savced51LU85iPzQ26Fk3kq61CeQ2/blKJk5NxaFJrd8nqaBqnA2QV7Gxg3Z07elc0mqw19R0bLn
B73P2qOwjT2AOHyO346seZGR0w7YPqWbphRhU+3yw3CJ/RFOqmU+K9zvwfjCg6HjRzOZWCoTrmxc
gu2/X8raNB3QuqRZFMFo+olMKBaSjl7nS4oIchREGE65UseogsMAImEgO9j7tCPPxH9cLS6NMZam
90xvI0kjxxmui4mKn/Soa1kyK46jQnmFXkKYe4mAE35KQgSFexqSHQpF4GlbZHewL9ywNTuGXvtS
oNxwKuByyfBNE+YPqdsUmuGhSBQ8Z9Fean1AkjY9zMjQuO1ThUpDE7pwuU1VhX+vgIRGq3/eGuLv
cDfUKOVaEgHOZXy1m3B8p6GVkc39z8WRbdoxu8QVljaHXeC6SrJJ8ggxBjoNanKIDTDOEIMyuFmt
0eXCZezUl73FHoiw9hsrSG67+avSkjZJvCOXHyNtRjip72SH1kRx8/qLwwmJDUDgRS48cLyIB8um
cv+mbrFSk+ZKWRnIOB4PqCIYKneNN/6b+IZpN6pNturMc9Nr9Wtgh9ZbbKNVuK2A8DdRdr33vM4Q
ffEKDnB1vYOX709SFPjAE1724b2zE5Cud9rAQ0vnBDdxtOkMjBqVpp01uk2GOUx56HsjNSXz7RG4
thieJxX1PVX26ZDgyAsT2uliHkQ9tritTqQbor0QuQZrP7uIyX6sWgLZJIhmPjD+n3vJko1o2sU6
V2mXr2K1ZGYMD4+wEr8VTcdHglzjNUMZPa04Qjct/jYfWJRrXK9LtYbz7tbnscR976Nf4Ck6iHJt
JS/7gSwf0mnOu5QZrP2AHlzyMpb5HU84Ly5WVJiIWw7zJ10IaoO+ucQf0FleFndsDVKnaAa9lz5N
ExPlbAjU9jJu7Z5yWh6JTJivFYwJ1F5ZSW/mbuEv2AGUgBuMnshRQku9T7qgqn1caxLcTqcuBToM
nZpV7rIsIej1bofGxfubS2NwL9Zyw1blUl+JKZT0jx9we35ijhsBhnWjpZ9oQD1R2nsoMFsZYNvH
5rCJvUkpe7lbvALt6WV2b6JKKrzF17HxTNMmjIG4IgXEgDSg0vJEl5ysDBCHNw1VRLOA3OKlEmzA
QXaxxSZymy51fE9eiD/TiSJc4LMKrbYHZoVL2Lyixw69WOq192lw90fXdUGBojxyH4KKl+wp7x8R
z/GNOwxnIhsSlhAXhG2pDguVkvJRYtB1ohjtwCc5KflSTsHOgUW9mu105Fyr+A3kiylCCfXBnw6s
WpbYYVR2ruxBNB1B9r6GLRFuvgunqGrjK58Pn5+0MU+FWgK74tpaYXo8pRyAyrCXLjl1nC222kO5
jCco8YUYqVuNK4DSF4PEArg0IME+Q7xTUVuCPY3iLWqdC6b0LsRPb0YU3cXCU7KsgXyqeYH01Dc8
yUXEAVujdMZ3+AHFsAjgkC3Mi7XiKS6wSnlIwzD9hOEQAgZS0apdVDmj1hLgNqRh4Jzlwvh3WrcO
L1j4krWSpOyO2xvViuxGfQDlx9sy1lq9kdZove7hXpj1clx0Cki0/pYmb0c+QEoipwYV9/f7HqDB
8ARwRC3wdATZmaDfAv2vQskEAH1Ldx069t2Su/UpqqygohuLTBIyzal7dHZKtK2zKjZ4ND3OVssM
s444sBL+yzA4fwsSXn9RENrPIyr6hs5r8dAR27aY0luX6lqr+pZomnO/ZICjMjBRAng9b3cO1PMu
85TLZtfLTE3/lu+juAhz0AXF7H+d/rZltinwR1E3SzB5fiQyBEWPyMrCJ4Hs5gLXqPs2opETdpMV
X8OLS6w6XasYxHDu6IBKggKQOEwVRgvWAKBqNtYvkRypyw3j+xU27doMnCuzv7Mv7hhV7J93Gz7E
a171Kip99i2lv5oZTK2Vr4hcyuUjL9+v9JrHje/hc/1Dl5/dqxcj6jNiE909eTRWGDUrHrXdO+7p
E9PR/lJ7kYe8nPjFqVKwN2zwCJ6hhnvZIr6yIEiYfrg3+bUOR6INDnoD4/NPBgFHs+ny2rb4erxD
n9Sjq5G22OErJcCc/Mq4Nia6dBD43578SMTaP4995jnxwazp6o6kkzMllvGxGNz63SJ0VFAXHStF
l+RWND5eTkjPBB3muZAOTr/T64VBsYC45SKWEnPbkeL6zb5g9DERPfIsfTO7FbG/YdikMjboMUfn
rXX8Js7dmhM0BFY+TR6N1Pcda91qdLbFdsmHda/Ei8nsxxV7B1YTwHC5h0hYOUx/qXwa2fEbQKNc
VFJkMFUYu5W0mXV/bt1VGaYjMTQ4pQxM2w03TGadIkBuL/E3pVDfbLWRFCTD07ldZm0eTWMRTRUo
mtY93Zs15YkDWP2OVwxPolzJvdAB3f8QcaIMG8dSVb3a9nYuefPrhX87H66M0EGJh41l5NcDwmIT
2yacgr1+laS0MbxL/7jEgpFVN5ddIUJLpij9SI7zRH2L9Vub9MhwTUk+LlcUsDAND2L1hE/hogXu
OycqW5UPKtQj2H4XA2q3HZo0hMp8l5ZVQgH2v3Q7Gp//cnz6VRBKCiTHT2qqR/jh8arcV1wcV+ZA
Fhd0xdfUi7ZkezO35UCBvmb++UCvINVgiJvkDQQj2w/ZYp0RBboVavcQtaNMNtmpO6KXOi374MEG
FNzP0KI0KDkeVoaP2QLFoaHzMHnkD3XdhOJlp2whUa0yelLx3GMjSJY0+7SyF7nlXBdC9cDfaKtX
SNKnC9WSNo9jbQlSD/k0i+8U2FVfWfIZTw5+1iRON2fwY1eL7kOZ+iLc7kdhjkMUOJ+X7DVCGFbB
VqNwDRj433ShR799KFtLg+1sbqXw9W733MeuMDbTbIajlDfo+VPglUwYMkLBdXhTLw6LrgYFSbaL
I3JVXYAAuMjF4YhJsyWhj86iqOjYoxKsZnBfF7XITW1KIRY614X8o+lU5U9t8W3/hwq54OGLbad/
rlYVQC0RiuQbQJCmIdbnFlGI13t1UgZrv5vvDhZ8OuxpYBXDmyPiAg3wMN65xRONw4dJCArArPM7
MdGedNvlbnCxo9FjSx6VFMyx7qYnNXLQPJIynjTTQhNnvFMswW6AD7DHe8NSZAXUwuPI2BYwjqwy
4Fc5xqU5klsnAanrl1KtgHzp2sfqYqhsRIaKSEngVRLFngKugEI+WzWf4Nkajmtdg1pRiToCF3dj
xtF//0VBm46GIwqe2anOyveNM6KRpblr1t4oMIAMasVM06DRcrVgFApIOWQ0MveMTuNSdn6GEJlj
C65wlnBC+dBgnfse0lXyciKyVqZbPj658CKmGVbFjZJs8t/eNecSMVqW+EPbzX+31GD7qVLxtVfE
BNgozyJWnL9oaCtNT14gXyn91LPlbhLRdH70hE9+FC0Jhm0QG+jsLQ7UCY3QApzDKg/dNEmHxK88
vZ3Q74oPrddRGHiSIQ9RRCYBJSxLELuP5v5nqARYJ72luZiO0TDjQlEmFTASxVkfHkPGZrf7qgzS
43SbeAFeSXLlg2FM5nVrj1+wHfb19VHIS/OzZVX9y9i4cKYxJkLWEl9uAYDHR3vCWk9H28FwSgga
3j3Hx9lBhowsZbWIHLsM63CbuVrw51S61OXl7Ro0HWzI2qLzy6KuP+uEYprPBGu7z0UCpBPAEieF
H4ABnEWV2wo9P/L+2ZFIcF0rPBGZjae6uJJ+eNnsOs9bCXn1veSlr+0IyruemMHv9/Izu8eNr9Eq
+k2XYZNBbNGoLGTiIqTYUx7nbkzKdLqO5pFhIv+epZuzfP0Ctsc6389CpgG6n+/ODi3pyHro7KxK
Scw4oGUcndaQSdRZ4jHkNbutwX2qRjVsOl0lYFVqRTlp/MozfMln83ynQLXXrzyEtjFLw9UliZFv
3/lRwKULhCOfaTVnYhObnrhhc2PyI3HP8h5zGbaVykp3NP4SuDGrlTYUnnILZZRYUUIrmvYLjGZd
BohxMctwyectT25hS8jOSap7mDg+DIiddAuKz34IXSmL4ZR+HHRs4I416ul84oVzsadj1S+QwkeK
jAT4fmOUs9By3fqTfsQWGT00Mbafr88XhIjxmRVuMo65ZtoyazW/e8AdZNmVvbmSYfTx/xUfiewp
EJRi2ezlHUaM7kN6E/tRWCItc0zDBfy5v9lWvFFAcDMnXhAHhFL5uiXgvGYpEfqCZz51ohlZaCWR
GZQ9W5A3asdYhsNdAS8wL4VEn8wQ3GZfSEmvfXFlTb0HA8O+vCTNav65H0NynUlHsAwU6DR5LQIX
04FAyt6rIRPJi+7WV7wH+uWPdSOjLWQ8JjW2fMYJEK/mcBSR4J1ak4VTCtZlYDQjPdpDyyBctWgg
ihKoY5MyVvG9l4xvEl9ReVChdqxko7vSdo0xsGVQaU/ZdQoUmE+E/0Vt3aygo0ngN2VIO95WSNHH
gAmy6R+1R9AsoLbL9UIdFaP8/vxrUFp54JxKYKBeDgfsscyFlgGQRCSewOLL2kylvIFj651FxroI
AlXEaZFNv0tFGmdihxqB2qQX27KlcSgfOHDDXdj1iVTC7ZrPp2L3+SJwawEFLTWP/k/HmYzFToKL
HytKD5llDsAfUd+nMWqJ2mrq/K0i79W4Wy9NJ1UiMAIhr2rUETI52fbHi+mX47fO+3vXtgFEdthn
4fuwSgdMct31+CU5B/tsSiPPL5TBCMVPfIulqMqbSUf2pdNvZgd/aZ2e7nRIfXtN5oR1ok/ETb2A
Y5NLsKdE3+pYVrEPr0ChWA48UitO0myrzIZFN6KkNpmmMfDxzvbwZe+oqZqERR0szh5uTW6/qMgD
JIfMZ7ok64jlE4VUUE5wHgS28sspODsy05xMI2ytflhXWV3VdZ+sJF7qF3N513BJ/KCDSLnZaWTC
fsQynoeSWah97jAHGBefpZUChjxGWgQwvoFp2Dv0U1WyKDui/M/WMJ/q1fs2iLSIXpSG6UHON9UG
1Q5UzD8tfUHAKBGtLgp/z9NvYtA1kWepO0+tvAVUcp4b2lOj6s8rZku5OSssEA3S5CV41MW63To8
mEALu98qK/XmehqGPW8Wg/Dv6B98XABdSMLIf+bL4yxTJNHPtHr+cJDl2st84NccjKOB2FnMlBSB
ayPf7FY7teya8zy8qZWSHbX33JgSSubK0egKbQxO8hLg2ywmpQOpCHaxrmm4+EKX9YI17wgannGG
FYE2Mnn2EAQipQe7BaLer5EePx9afwqcONHOUi0T05ohvnIyKl0HM3ZQCV03Pzf4GLcm09BetZAQ
XEw3QAxqMTP1oeeITaUTaaiO2ZgkOszvoeKQX7dOrAaI+RJhLAHbKrjoT78qtAEFBIo6I3csmfmp
VZp7DOiTPBC7GxkVdd1FuyiyautmYo6ndkIxqqO2WK+4ArwH1bxfn3P0TVlEr+7zaEvFKHvOUvnC
lKuqWihA1w6TlOw59794btsx0iRZnR95bu6e2p/RSlJK4CQUC0TziEK+tWrMddPcdXvLtAVxRRVF
/4X6QFHw4S+2/EryUWPIBtCO1pqW1REJaM1W88em+rOHOsStejyBKb1cl5gr50LceGQFBvTCwJXV
hvedjtnoWKXXPGgnW6uGxVdzSMWSpjeDhV9xhQsADwHCXcQOXQgF9fG3/WG1WBe4nNvF23x3CWjk
DYf4LCGDSmFzgclWuWbMILXacGQibxSe50Godvd+qbfdYMb9MF3yVKk40UJmRPJgATCusFQ6wWWk
n7jAZybeQoIAP98YtIeaBDR68KG53fv8jBwGRZ5Cj1DvcMQr0FkCVWzHL0IpFkan3ZXdG1ktaXps
+vs4L+ReQgEQceP71PKZLxjfWISwI3D4mpocMtn1tLXzFropeO32McdvEgBvIdsiYESxI8r5ZGBy
Q1DDz3VR8I2Z+yjNr8Nn3xWt+aExTeOFHNweovjq3ks92cY3Da4U1btZdheDEwd+7TDX1RacXSgp
8j8ttbq/0uhfze0zWmePEmd5rpsB+OeEiB2f9tGs8HgDbaF9+OQHOrlsndjN6Ea1XfENECGepE8R
Q0s+zkilJkv5n2CVERGeui4kA4HtRtGIuU/BrQR8907dfHTgzJAy9mOw6v3OGmd8TvnlQ5ifWjPO
Me1Ld/hbgpcct+C27HnBMNDUkcJRIQa3rAR3vykXzHqx9vXjxDMF9qDKaSpvi15rqkx9e0w2ZfgF
AC5lptTWPX84E5wz2JK4nCBp1osQwWfV8N5HhgH90/APY0FkvpC7UmxtlRZdt7R3ex00eQtZqX6X
Nrmyj7Gn+C+iWxMKSik4fhYrXs2TcEZ+rAqZG79ho2bujhRnA6e+7iSOGuFdA6B7nyTkTq7BT64i
X03+tj/nUx0xuizY9OZGL/G0/V4jEIjzdgqlrN8KPi+iCTvNNMNrFWoPO2FTlVQLT/WR4fXkM3lT
fKAbCknzp/yaPiLZyjgA8qoSLQrdGgKUdoISU5VpDU0MUHXrMS/UeEfGIuj++yMObnb+pouIIq+n
s++RrZOEF+312KVnSMiJfzp2N4ezFVn5SnQWWKutHWB3k+9yHa3ciWn4EVgLyaTPQ+4YFtdUlA2q
5ZmPkClUf0wlkXy1INcFFtM1wfdqN30MLOBGOlH6hd3aMcZfy1f12GoN51SjrXpnPBsLin218PIC
K4YXouVF64VPrqXOyG0EI+jz0Da/3Xqb+MS+UildV3jHCuWTY0pA8C0gv/00vo17bsjuEN9BRNJT
OGiYvX/UQug8FOFjRW4rKyln69jwuvcykdcjVSjZyORtVdDiY3gbd+HYmL7ZuzvJkYCPf06uclnm
mxY4XGciDrlngNaxPuK7uTboP73i+OCLZh1TCCTAPqGctPOIvbe+WDFIHepR4NpdCNQwrDGY2++3
yOMraRAgmU29EI7OZz5YOT6DT+OM5tfsWf+C7w4uhj4FkuYLbZg+YJ+Plgwc43VPf+GXHhZ1plZl
FlrC8w5hw2TXO0HUCo2B+k0/WlgkKDzcqvc7ybRFw7KPvnvS39qRNnFI33Deu9VTaqTEthRVoGE6
bQt5k3tBYmfL2Qwnqd0ZSqdCIC3Q/LABZemoj6Mv+tNMQzIBzdpBQe43TsXKNCpBKsR+98DmZNfj
NsG+j3wXJzsqpbOYBQzH6X14sOtnJQJM1h4LsZ0F78wOqqBmCPjEeJaRNo9mJyU41pGDC6cG8mNU
Ouwub0b4opvla9QIZb1PJEH/Z7nuzKAQyGEF32P2Rk4PtWbBJ5KZsfP7Yguh7LXrf78VUvwy0phJ
BRJ5EQ/jKvrw3tD9vodTL87WQL/njzEkRepymOCVJSpTLN7amiKbaZf3ZRJCO+00UX78dpA3iirY
c/i3Ng0AIUR3yM95MHCcv0eZiys4K8pWu8f7YMvr9tvg3ac2lydtP5GMmvtIEsG7l+iniMsCPUF+
Fw/xJOzIWFQJN15qbpxFXlXjKVqY3sVCCmDACyyB431s966FDPTHFliNTJvc0x8CakrJXPZVr904
Ht0Z7bQetMOHkg5jWEVHx4LGWOL9oajHIGEBkuArRY0PnMuqxejZys42DtMbyIW13TWf5IxbmmFd
D1s5wLM45iO4ttOPJ0gwGsNcBh5iNLGG/GbFnLtRvQfkv5mUnNnxPBpSCzFTiYcONC7zywLztUAO
Isd9Vkh3hQurmDTSMpbp4UvOy18menHYJYwr9DtTke/m4I+gGFjR2xZ1Xj8qaVojZSQxcdfZLJuS
OLb5iRs8PZGf/vw6zx2d2UaKjSywX3DD423HKSuXaXsCblIPu5pAVRT314iESYBuh+Nmmm/kSqxv
8GD/shgF/IsiG8TdPq6fTPpnEVajNd274uoZ29qn4EMOqgF5kkyOOUaqr9WyABxvquFbDYpPnv6O
fFrtyQGFdzkbbMa/MXXhqEeZYXmfle8wlrPkIIAwG4yU2i5Xft9vkCjaUaQL8+sHhMjTxjmf7c2l
a8gf9race5FumIsqp8VLUYCGHIZ3PSx4fBXPf+MMQOf5mEtbrhdjcgwYLFtzXLhFBbgwlYMUwNW5
HmtWgdDKW6FLuhIoRv18twehKzMvcXnyEM6hIJv4ZiwjWVM4hi7wXbHTMmJZAdR4Lxr4qx2UMWom
vnSht4VkWEoZtRlF6tolY99zSlOPc5utQ0Nnn85MN2ixta9tPHg0+eAyq7dO32aEyXBIQKpz90/2
mboDD9L4LWVx7bM5zLQFN3eLK12DyOmK+MLCVuZFonPrjEOi482hVdBILCZreiW808UIT2mRVp9o
k/Jvb5vtA3Kb7qgcaKJ+eKkihhyCGWDTm4g1XAmJFsI3PTBYsaRwRTF5WIIja8uFJuTOodY3JZkW
HKmnurxn6CoG6c1U3oMyYI0MYI+1Ht/ZjAXq2fTpyaxYz5hBQg0Z9idwFAlnnYKfG2h6JpYh5XCJ
z67O3EnUvG9MkBk+ivxsv3at9FEJ9TVTZWufpGdyjdIdGTco57DyOXgK3fBTF/IqeSaCe10G5WGq
ctyOhRsLxXcR3vsKndLjpFONc+Yhv3xXT/8vfHPjLgYcbf1LgWS6Ia1hfACiXsj5zUDRqQFKyI2x
RhVwx/NV1vkxtTPb4IX0qGa5nRiWEs8NitY7A6j2eWzIRAgxTOe2uwelDM7GsXNhbe1Zg7VMl8yg
T4rabVQ1WK97N1kE7mAxanX4C8/bmI+vsyfViXuFtLsob4xSnFXe7t0z2LS/Xjeepu/ZcusKD+0g
5i/L19J0aBjC4cJLe5oV67WL0Xjt8+3OaWnjQdRCewnZyzOWMNZlY7SQlg/KlBzDlgZM+jKbVR7y
KeDhiRuQ0veRlqNogJpP3/sY/5SUyrN0lzugmVSMR9Z0rb+4Lq6wN70NoPgRkeoyhDDpAhTyQ752
sPQI2oKfc6r7hA+ZVXs7d3nItkLBhJRjfUTLyKomUaKygboPJXcjshmWcuE+RuzrAtKo7nVhEJUY
xYfRzJIabOGNmG3ieCtM2g0NnEXNNqsZI4lRpUulflnrlKlVflF50UjN8s4fdgWkVQajnPH2bL+b
Z1dq+u7kiF1VuSKLYl8egLZK6LZdeX9EqqSnOBlc9pjQzOmJCdxHi8IK46DPJ9kMzzjx28SQ0FHf
42W8E9gz27ZGl9x3cbUARTBQgusymfRUna6xr0+LX7VSx5LvxHPfegpwCL3ZMozkTMoRTb+op5jf
0Ew3K7I+CI8iEDb/YD8Pm9HXB8WEsPfHKGoJLn0quVl+alU2Mdc2Fpx+y4PZhIbbTrYSNaB6+4ra
qfJNhopIXQYbuLfHKtqGoLNSLgxR3nGFMpRhPzSYManJU9w6tPuuu0xMRMdUL2N6SE+PyMu7na5D
vZGJDpuIPaKuDZQWcsnn1g4XatVW045vOo7QtQ8L1fwc5k5YBD3kZO4r9nvatFFVllcYJOMRTQyk
NP3Z6JwfDy0zLPG9a3Nz6kliQpq2X5GkT5+hk5jegs3DTeljuWVjsCxl/m+0xxdt87K3tYRmwWtP
JlP5Vtj+KpKhD3yO1k96puYvObMzCS4S9ZuFgVr+h4yevsgJZjzqrt3dUR6FNny6JuD4WMrxgSmW
0zOkSIk2DrcXRJuept0GrR6UKIu02vgPftugkrD1PI3bLkRHNtMv2lKDm1cSDHJAUBhFOQoHSl17
3SSvo9IwkgxknZ3NtmQX+BD9fXhKtHV/scHhvjB7WeSLYI1B/eAMEo6ElJOygqFaLH+aybU87ZXx
b6gikK/tK6MkuTLFQX9BojXp5z97uv/IJRgoMtGYAADAdDVEPTrh3EmipeKTFSHG/8tZu+T0DqKE
pp7I1+PO0iLyIkvN5U/8GUtSN5oDYgAOe5MxNkQLy8LSy848e7IOKFGgojE2gIrUvSdlEj7scmnp
XN8d+vyBuSc02NiY5JDArhE4SU1MH57DqMwCsO+Bfad+mR3ZhkvhWnqVVi1jZG05VA/MLAyh0YqH
J+XlObVoic0mJfZ6DKqdyqenAb+XBt8Dl6EZ5cjjg/8Zmo/m8pTXa/l5HdmvwVScYj5GabNpumwP
mw2oVV0ujbXwFoxfjvHqK0DVJjcNOmupEGi483/PzdQdjLlQuKviaLjp7ctx4xPgejp4AMasId1u
rbjhbzyaHd/xVVgrQA+KBgABjqZyuYXqXTeJiKmAVSJ+CrqHRVLcBybyk428qXAsOD+aQWfj4V+V
lFpqEHZEMDgrJf7lA/QLN4iA0QRX90OXGvmb67Zqc//Ggv8/MYD7RtrDuQvw2r7ZuqR/qHFnuIhu
QPmHRL25CAKbEO0NWKfMmGuD5dANP4Nn0lPg6UrGVKSWpZHgoWfEWrEguCAhSRXkIJo0Xh8ctQIQ
4u21c+dh+b0ypbLJ1rng53dKyAhp6CtBL5z7jspDLMBSuWsjScex4LQt+iVibuiaCma2j2EhRcmw
sWtrQ7JbfynBNSwe6VEkohnhrcVlA0x/M2Wv4r7j/LmUZ4UN+ZNpZnp3LIwO3bcbnIPBPFqQK8NZ
02imWONkMaX/Pht/Td5m5vdbLq3P5R4kOB2AtC7AN+jJysvML0mnoqp3dem/TGCctNk0Qvua9B9I
IwRcur0CNmSTmP6VbU/23XAoyKM80E6/CK7vNt0VbUL7gcV2sTGO5sKtvyDIJlaeSi/vuoAAsiTd
LRKLZxNd9saFBYKLI3mVz8ZKyueOIkbfnT7H33pyiguzeAOzBcm9+dWybqUezRKW7muLQw6PtTcX
/JzpSyyigDsXTKqqR3/EPlJomSlPQCk3j9YUyl4bpPVTV4R5uK4hIa3I/A6gdyOXMcyGL1gUISNC
UTG+GZbo21IbNrNsh+FfKJ7BT6iKApCUxMY22IjG5xcDQKKv+FD4lM/fAXhkPrN8F4O93TbqP29X
WwafFZDPb+02vjOGc0f4eaFBsoGUZfyDSjFzfjfl7KPog+8VUKah6HxRFyTOBLRV0tq215KZr/4u
g+GKfQpQKKDOPo+QxQl1SECgttC4RnizUPDhrCH+3gf/2gBXlxldlp3G7Wk+F09bT6S/kZSfCY2F
Pis2wdUIw7uUU5R79bGsktjIslZ+hYYE0MTU3L8tW2enNsluvJXQhKJnXMaFNzv4Xc2jG5axVdGE
ZT97PUCU5rpM9Y/u0wNxJDySuU++2nR3maIrdWBL5L20wIy5K/tagaWNYtEFtRmB85Yg9kTyoz1/
W9xM8bpKjwUUXYfoCczFKBJTtDfT5QpPShd/DifSpUoqeUBQOjycVlkjtl3AmjAN+QTlfXHQaEcI
sbZ+KvOIvQl/n2js4sMTDzWqf8aOpmGXCi9scPhaNwpAneanFHB1if/xA7j30THw7Lovo+aQrn5A
pXYI3Ion/k004g51e3Q0cEtHZHjgy2gnSUlD4mJwUB1K9z0r0/QA+mnuDeLWUypXMw9JyBFgskkn
QDT3BonHg/Hz4YSPZeJFztlDChL1XnqmftMB0Kq/38Y4OyjCUixtPVXK46AWAUplZUCiR7vB41GU
TBj1nQpBCn8kcCk90UXeC49d7ZUOTogqi4ll5PV+9YQxZM0pmheP/an0Eiw+GficJv1P37KVBf7e
qdNI74V83K3L0JQFD44N39Dlh5aC3/C2JVNwVOfPCeQ/EQY0J98uEWNZZZa5T5FskKL9ZQwLpRh+
Q2Rvs+j1aW8WNRf7teMNPushqr+ho3zor0yiTznTPU0f4ww9grSIvvlKLRuw0eBN3L0vVr/Ymu42
/bNH7R/w1RbbVIKf1zRQt0hDGv6kpw0XvmTBCVbbKjirxOsqaDynRf0GtAsjdtODxmy107APpWN4
roid6ZnlXCBKerVJhmfD+omKb8JZplOMKikdS5QYZwHPTIiSMcbrIuuDu2+BUUF6aWnXJlh2Qe4q
TcJ+hGRW6uKEWBL/OweG68cA6fXuwvSXZGYn7SqonKIr6mM3V9gv0o3fXdpnPjjuqx+XdQjDL57n
6NFO2NOFXda1XbLic3by3qBA0uz0nBRdSgJx0EXdTT8QjgEKCNMj4RQR1EiOUdUgsQV7CMhw1pFT
3W0g1+n5fhfy6IVmcYu39m0txhSRjPqNNFcRP+q6gwAxSCLV1KfpWGlveTp13NiBzZJgY9Uas3+o
BXLXN9EIGktzVzMw27fMHJzxZ2d5iLmRoPz+1LG/Ww7FUfSXm5hO4tC3RnvX8/z5pl8ypHfTGOMw
RN29fN2cwNDh3sk36wCeIgeF3qVSkahcKdFgzzl5IC25lEfl/GIGgpOuWx0+SdpNIb8sNLs7St2K
vPNtehoVA0/GLB6jFS+CkfyUrJwG3j3QBdj2UlWAYZxMPFpReIO88/xt8FXwh6JI2cyxlov4YVT8
UsMysu65Wc+CT9sOQe3TgeiwF+ORbxWAUXQEfw0z7d/8ccz0evl5Wu0HXRdzNyrRQdQQ+LkTE2Mr
6+YsodttG4wM1AeP5W7VEl/8+RVr4rp/qeD0Zui6+btCqPXx67s0KyzG9p1JvcQHx4qF2PKuQDX1
EQhsiV1/vZxARTpeT6KMRUq/86jVaqNW44PEL5wMRjrwdDDGT2lG+n9bpYTtm3j/G2LL+F+lxUT+
icF7RkanAChySp3di3agWZiINCYVsymFS3dp7YIg7tpWyls5lDDcY6JyKE0GlLrnBWr97FMBhN08
Ker0NyDQKEhfLRmhoopzhTyq9FfVj+O4bwbwZUNQ6cOUsIhkQsM7M2XIHpXd3ZnEVDy0VFQZ8pH+
HIuTqnKkzbP+OGacolXAUmMrWso+3+TYfIzqCbkNjCYwlOJJb78UQ/noVNmKseKeYYNZOC4YGEbW
yKjs2WIdBa/C30cZ9J0y5eYQreMGEqu1cGNOptCTFQ1Zikl5bezbl4zFHECEdVRNhAWVNas6tIqP
WbaPQ8awvA2tSCRSfBIoPFlprJD7zF3/Ayhl0gkopjfZ8YN1sz/7YS4HN2//l7PuCHB7r7yQ54D2
Yo5OjBN8hkHbSjhEG8pyUNP3Wrd+kuEBwjknUo++UyNnwLx1iyRy8OwalQkYQb6tzFfFD2VqUbMm
YFeb45z5dqjXrvNzC3Az0yBWjlJ47nlpg9BeTg9Nc0n0cfGKDrWIROA2EWLp7yID6tnZD1Zt0lAV
smzgblpvq9tTr2gMUZu4t1Jmx1S0fS+UoZYe/VpzCxkUEYiKI/mAoLSoVK55L5UAQ496O9PrblWr
cadsA+OWipv5mVG+ViMwOgZWhK++y5B1NkfdyBDYQgbBHAoeWPhRBovPnG1IEwYAmxKFcoqWDoTY
34MhdDGFfuDlKNBVOb9OPM5Mbw5szD7zvPeOiwr9trN2wii22H+K5AYG9MiuurUl6kf7DVZiKnR8
MhGbPo3ssGMuwSYwj1k7U6Y74dIOMno03qsD69dpb6DNffnGLQllkxDSQtE/sPDvzlPwFn29FZyg
rG+F8GixePg1hhmJATOdXHp+PahMDzqUnnxwQQHImKT3EFlcw9ibgQ9acFazPBxZ/xZZQoD17OmW
HKwr1Pv2Dgonf/h21YYFopugW3VkmGEUVuUL4oPe2QGAiCmMQuHfeX9xkxCDH9uRQ1AQ6e0ceryn
tHI+RhAW0ZTx5/5UC3Aj4SBpaQjYdQ1+YD/mWwBUA5Llylp1PH8yTWLeF2Nig7w8H1nrnYOWqY6d
H5bLi8HMQR6EsXFsfDQOqpJ6r5qWnImc7q8J0cCNhy/fUKFmtFmmEG8nkeuweL10Pxw/WVp3vc4s
F7NcNH6E7IKO5P9gPgze9nFUg6weHNJMQ0GubMq34pW5zO91Zy5r8lTOgkRJrUaw2FofYl3Pz7W9
xTHsXcz3Z2N0p5YQCSH2ug9+FhPddxVCxWzMBGt/bmnDLY5bf2eKhl4/DKSbhaLdbOts7zd8uSS6
rjE3nXMgl/cgejFwL+fA34E0a22N2KSNadRHGTuayZS7GPc85+E5z4ZeD8UkZX+ndg0/w1F+aG0F
hAKqC/pCZO5ABwzvlqBWhlf7u5oEHdivs0ikC6qp1BK9Lvi9bqcJAuDJe+nQwPWCZjARsjCGAS23
ZABwKiLsOzsPpon1C9cvQSMFsRfGMGxG7gsKVtLVEpjqHYrMQAY+GbvDT6ASsDSIOfkgHn0gSi9Z
QfhxxRb6ArOFHDGi5fjFrtB2RJ1GvP6KjwusU25rpIctVTvwg9nVt+2qcDq/hEBBz2wu3QRQ+ZFS
kU1QGS/stSSMauRC4Kiq/3iJiUDBeSnSxJ1SxLVGW8VTYvYRC4lpsE4gbbbVQqu/4Zpe5F3JhGaw
ek9WhxV43pFMkxI+SZvhFnDEQfCxHmUCJ7w5cOTX5dyWOqAp/pRpYg8Gdv7zyZDqFt39AZBlC/7t
KN6pXwnp71FKrVGtv/eOK6A+4T8z/D7X4DbljCnI/YqjNJ/jxEWzZuPOy8VKyWohuEppAFe19irf
f4hkywP0ZmLgAAVWETk0LM5cAsh1wgJGE61QXS9k6X1DmAIM2Lwa8BET+Mb0anSnjAci9NLyfkUP
7T5g7hEOqWBRvNSR8WW069iTT5oD24hyWOlTzvUq7cCpckvvYSRzxTJ9vK2eochnoCjpAqG0MNrN
lTk4rL1VImwhp97u5Sif+If2o2Nzt+oPB/CmVWmzAzoE9ioOcva9rYXGeJAVFrZNKksOfCE6ZiPt
+tXgEg5zNTX8a24G/7L67yX0ZY9SYlBKBWrtEr6LqOeYWvGZXwd3MFyy1o4GXMyTrEmea9++efKD
OkaoMEMTw/n2exS9VH1MpGZFx8jugFk7VCBkKbXEaHrugqYelNsM3dzi0IQTxSZrtAG1zzW6JW6N
oX0IplAKAKHFnQgYBc2ZWhotnmoB6NZQzFuDOaIIpxAuQRACRqGhCRSkZXzbJgX3t+jDUV2yYcSC
bgWJHRstUk92KP4HmkNwO0GBe73jDpEsbCuq1qondwty9WWEyMfpeoteBUGg03ZOkDiVdDQTHx+6
BTpfPTxExQFpS5wBVAY99FiwDv0aUBGOTJbMS8cDcJPWYenx+5pbo/mw0rrVlamKJ1X421C20+2N
nA9YfbNbSALDR6mjTGoHSBj9cZ5Nc12lI9KX1lLPi6Bh6Ix7ElEEHd2EbU+JviBQA1z/5ke9Q881
w0WG6jsLfd7c0Jz0K9XVudZoOBoTbIyiDoM0c74Hh1Qfzos56DKLcm5qD4Un+5uZwyLW97aX+pF3
CAIIhobSE2ZAN7IgAU3NgMCwyHgi+mzibyMefB3FIYdF4itETAkPiWiWqWULEtfJ0F0vRMX0SKhQ
kU9qGP4srupZtflaIUnPC4IQ16BrTPmxBFXTg/aKN9jRMt8lR/pSbY12Qzym6539MNcQTwHoAyyw
NywEHWC6JCAjr18YnoXEnu5d1QTLwnXPf1LKWC1d7rTtgG52maC+TiPMIjPlamD3shZVm47u9Sh0
Jm0GAMpguTcLyRfhlJAXmDs1wugbOT3hGPqbwCB4LFFdpg5WzcXL0inycnz3eGFZOaWrDZ8Q3jyM
BEyZyfi2rMfQTStwhu370WtsWeRodVHeGU3wrH1vKTjPKpj5BY5lREWmhIkFhsGpbbdRNjYGMkU1
OyJdlyem9yrvf3PyNYbpshGwoU7bmaOGRdtKzbJGzWWA9LgdOTaYEVNYTNNkNMxhCvgl24RLFMc+
2FtcU1u3SyqXb1yUC96J8wYzA6zPokBThXmFZG/aDxz6Eew/XnFNx6ITydGHz8Fk9JseEICdgjwo
rGf/QkKiyLv8hqgmfBplOw33YzGuETasYrGzqLBdO1M1YZct0gygZs41HsNw81EITZnlwyDcXLRO
Rd6P27oAzsmguyOEmD79LRcf1EPMm9KK4ggjBkQcVFnnUsZ3LQpCua48x7l5lOL+9egDPaIivaag
BRzFi0h2Jk5txmlfbPTI2m21RoTvVWDnGKUDetvA+8BvuP6LaKovDWHVSUzMVZKKkoUYxb5EROZH
NSH67Wrz9LDHzxBRm9b7FQRs7P5ZD4qkIRLRcjb1gheiHJbwMMD/uPe0EMG6Ac0MfLM+jW6fx3M4
nu+Noo8rKRwOKe9hL1O+oOYXzQntHwTIlaGfesmIdrIDT4Rggg7JoSMkUj079ATJZTtkylJDaaHq
TlTnjqWeVVTILDNAkGJGuxnZYTEUR2hmuEcUzHP9XgnlCYpEW+8mjMQPTrbCEbJ1fgjwGj5ZlWDH
gkkJnkkJWaSr6fdhmCkCALAUEqgNTdL6SH5mEM6df/KOh4V28wsgFHURsiFQ1hGOfAaCqPNl2fFd
35zcjscVJH0oECYgkB2gnIcGbeUQyzZc1GDzw1QnuXiuiCsGLZhPhwKKdz93DbfbXLhFsNh8otDM
9G3bFsnffZr5aNT1MgrQlABotU9+cNOiF4nTH7Rm2DhKlZ4rS/nEukZcufMvgkxpuHpf+DUJGQeF
23W1thEykBl+Dn21QGDRlZMRIFQu7X8tGspAmILfcGZ35xtGHr8RMNjRXSNEbtSO97Jbr5ml/cxF
NZKM4rGFRPyTGvpulaTQX1GIN6RaioOUkkPIXde025aLs9Y6OuFL012IgQCRiuSWUsRJ4Y+ivYHe
4rIB8R2i9a9zCiXiYGKee/W2W1d7fvuALjKDIKba1cOI/fTn6NUrAlyUMeB//LI5wHtadeWIAZlZ
nOVGI3jOLtPR2GsrSP9tFk+Zwwvc4uxf6I0L9m2YvkfvUFlgtPxlx/mG7+cLQmf2ypWJBKZUtNWR
g6ET2BjWgb7DjCJ+8rMrN8xZrAliUbzu0RbRoRgMBK1pkxZD1ylNMozM+A8L2cKn/+pswsJOqwSJ
XWqsl/oh1hAC5h8zmYRdv2tKUU1zZQ8OED+x3jWQbiIq+q/vmw8A+WSXK5AuCXOLQ9aYCRKiP+JB
XfaEQtqMfIoMXM1uNwHbWDSNKJRIZr+HCpPa2bjYnpIi9LAv9rkIa6zbAhv1wB6Ppg38IgzWPUrx
giBH3YJXBANYCbxfNBQQzavv9H1YRdmtWIDB495PsDQVJwJpC/xHKmW8FPS/rCuwN3qtTM0mOR6s
UKU5avigjcgIWG3gfs7omFlScsiLWlHYjEcs0PoeZDB/Ev+7I3AJtsswBM0mIqTgSiXidFqDizk9
V9dG2VU7qp4kCpHrri/3vOTiYqFr9oipGdjRQXaANHvc4b4QHVNMV8mPKBGzjbKsQ09Z2dJt1NwQ
iyV9ig4lMv2RzMugY6Hi1cEa8p8m+ZqNKA7BWzO56ID8RcELIvstdsdDcMja/f+ZhLnBYlaWg4fN
Kxats/uMZoAwWb3449aSZWkONAHhXB3K80ZosGnIcvrjtFQcEo+zHitAVYAv6cT3Ugo2187z2GQf
ghJXUThdSnj9LSVLJwAu0449Gb1AbtWJJrpKrm4zW7YiQ6TrrqY/KTQc9VbSD7QHePOiGupCDsx3
DAjEG/Nd2QjSOjb5YBhn51WOPAwub4yU0bjFEB6y2id6rl+HD/ltVD2P9SdF0D8YhPqkJCfVsZE/
5buBqCcuKuiN5WMI5AirlqXqCfdHs/DL4wcEgM4x70uDnLg08mzFek09adnBvfa/6Wh7nw2SYD/b
OpVnAnFijTSklOTxCHxR7T8PfkYO01jSLfeUJ+g3Ydq+VDCGglwmjA03pefCek5XUWGZAhuzPNOD
kEwJbhTcm5RQXOi7SQj9Ic28siI5HZQRKG16smELH9L+7M5fMw49nwwM5H7Je5Y6DnKfqf+Lu6lw
BoKH2fVeE3xdhT01LpCGefjmOgj5Z0E9W7e/WAjRwK91Pn18Iba9s9/n6qdopS8Bdh2CFDPiuBaE
eDKf00/1+bFibgh2DVN0yx8MOmw628a6GaEcWe7oy2BuCkGsBSeVY8wh4LfJMt8Kr23PMBZlLqgv
zutGpzYra+JIwX/CGXJ/yRF5S9SpAoLQim4e0E8Gwvyb5WuA0CDRMOt3G4pK/wFR6OMCrbdAoa7i
gRoor1Gua3CWVe1nbnY44uOEFVjeDEcZ0h24DmlWwzL/PVc+bdLkLLA7/uLgvqyloyDW7TVUjSgm
8Yel2jEGYY67OKprThCUOoAUG3gxDSA5suBtgoi60gjfK6AYhEse5WL45e14oL57+85e/Jc16fHl
Sl+njmlVeBHRw0tOYmCZbjB4IRsVgrvL3DlwcvsIfvABDblPGaWxKPfwjQM0k2dykvKRBZdZmOxS
bT95k29usyNANxMyC7WnIVMta7Lz/QX6vg5z6spv+eKviwdm1NaronEQhD9KMPwGGQnrmTB/VA0t
oT7G6dPNqiPP43WWtloLAmSSZ12Ovh7hAD/LCgDsP0GynLXgF6FJI+KQVVoSIOioTdKQIKiG3Ib9
kob0EQbVgKKVwYiWAglx8qHzLtT7XXwvdODy2ePQ0lWHcA/UH47bs3TKci+yb27osQd0nORYjU6W
o/Vp69A8cHNGoG74Gef8ARTKmlRVkMm5/jxhOAFERbxwCAaNHekw+oR3pFfnO73pXZfzPoBhC2yT
+bvomtedY7JDYN5IfeNuhGSQ6oKl81R84gyWIpjfQLIwBrin54p3KJEUjwuD0L1SGn8nnGZvVcBg
5OjYapd2ZG/aaxRl5oNjcMdDHUECVEIYvTUdGSzWZWB/gpV1AF6c50r6q5eHHUEc0GpKPrte5fvl
sI/oV5U3UGBX/fyk8i3XgGutGsNrAGShXd52o1a+DUh5Sozv43qk4UqbY3ArDSgWM0UE6+V0/wm+
qWVNCj7LyVGSM4ES7C3jirvwVWdC3goxZGtfQG89iYoCWcDnrlLBidcB3ZCgI+dDpU1togmwXncW
dTJw1u3qSt4fpiGcq4WVZDNLuJNtlNCLZ9CkVV7YZvTRZnhL/BM4cfDX1MzV4Llouv+9/hO/8HPb
6RGAtSaCNMdRxJONlyrmg+ry3OyGUoEb88dHde7rYMgZIBPD76FkI5Q2vkj/iEUdnO//JuwgrUw9
/sXAChwtsSScgnbvViIiF79hcYFUr3wXfuJDVVKJd0uHferzlBGDnNEYNbR5Y66xFi0q8B85fo7/
hSLJOmgAb/tyA3fyC3aAjvq6S6otSiO7Wg9nWOSNoo4ypBCU8CKo9rvz21B9gm8+Nf5NuoaquFp+
efTBdhpWIwZHlBM0aXBStFK6Dfi7sQEcGaXCB7kV2eQ6CfpP5AaPScocDmhjbUMblTxoW+Zc7GTU
57QnQWEyuW6ODzbmrsBIkJkJKawq9srsJQGvskaYoxzRevuGVjDLr4wxp/SJC1uvSVEBCwmbnNxk
BxDte0NJhWNLi0GEjA4+Szq9317Cc9EBjsF/AnO36dZ0XrJ0l/4YLjwNfhZQ/+/HerDNhLjCPYHy
LqTnw4bf/9qTdTPPSfpjpvmHjyz3AZ5PAahApITZvjQRTzAtXlfDyeAgjwGDbSkW/MT4bmJxmdd8
cE/I9O1r3H0jfdNgWeO+n/otmfiaSq1tUhzxQtfkzMxcn5ocv5Vz+B+nxkdHup2g5G+s5h6IXeBp
YP/mOK2rlaKzlkjK+jFruYsW0+DoBMpt81GmaLlCUrII49IDBoJaSIpeTWYnAjCQPqQvZ3EgDr9J
ODC+1c/axI7P8rk8W9+D8lof5rQPLyHWvmP/5fNy+lDHRC/n1zdcmkOaM9N/b8l5s6+P50oRCPPU
pvELP2KoDAr/qo+lo3w/Pk24adPpW/rD9fSo8AA3I9xOGT3jt1Cx5gAdDkUTiJ5R0knjBiem/22A
Ow2jBieJPJcVJupHcMV54GIDZQPMkfzroQVQA8xjdLQ8iF9n6Bwx+sHRXNhMft27lERogCic4Liu
P2czT6gCRTCL2hraQvGH7Di4KQ0mxRH77nAneh2NFbaA88d9f5SoZVLiPpRq24ZaeV0cPLcT7Jhe
owqcStJ0tguA63q3c6B6bTtJhWYiDwJPIQBzwh8HgJOG7RDpsYSAHNxUlOjhihrgUjj+QmrHiu3o
6XIQS7fsfqVpLotgifJ23Zq03hYuH6exp2rFL8pkolKLGKSY9IAuBfaaWdz89VbZJKTrrdyY5gOu
Q5TlhQ4GsP+sza1WPbD43OUxHkP/U0Ig4NVFyX6mxlDYhuSt8gr+5O2pblV/yihxunkrr4LiRn5z
T09NBtLCCYoy4LQ4sXEeb5ZG3RfohwIKzVqIEwQ4f6R29KbCH6BzddKhadxMNr+rsoMAExCfzI5J
VvLnrDaf80JYSY++NiintUpsRuSDnZK9EcHv5u6cbZxQzKUiqmTJqzo1xUQYt2mc49EIV4bpQYxx
6RLkl31BJNlG1Osz90IvpjnxgtAUPtPfDCiikCFJViVq6V0dWmaKEbR0JI6R6wI+NywOMuFkR1co
IGicyWlRCfOo4xOJjnObrNkuMkB6AVkfO2hVY7A9Y03ZclOBwNTzkGEBYkduoZq/fxbn/OebGyoB
g4Ik/+2SbjgmHO7fwxaK1QYvL2HJNMwCtX59k/cX141Zyygb9/a49Ic5FDUQAqPosbWF6+KqmCNN
Ef4Q9KClboBF6+XMvYGitsQI6WszR8vRMPGgc53GfgSBUHVS87RMqStXAs6SaiKwWCZzJY/GYqoD
AOpnvVLCRnjGMKDftBNaSMlWrtNBZbXt2epEninpoyCDTbs3tvveEHis3bGSL8Di95OsbfQTgbZQ
FxvhaL5BKMRGo8nwJHrIpwoshO9h8CRD5WEumkmU2HOHUbRvWioXUXDGRLV/LnGECV4Z/7Jr/CX/
0X8Tlnj9SNruo0+2N7yaLwPSVRHZ/Te/vhvO1ZumB4RqY6F0sqXGsUbv4nbJSuLvvMNRbb2vD8Qj
z5B7tnlWoL/yGo/G/26MtNj04eoX7dU/d+1em2pWI15U4MAWKeA++/A4js8pN/EN/6t36UWf3abu
4LD4qtIbpe5oHO7aSFmibVnAaD/NH0PkT7kXsem0M5HQbLPjfEyZ13ZKlVS+piDUiZ3rC0A4ms/u
VxKv0/TWl8wocs6IMjuWCicxlI5F9p3IyYtsSzj0xQ38mFDBMq7VfN8JHZBcK6g09ECu2MXoUgGe
dtbGTUDHcQakNGWp4qZ3RRIoc/bVotd+YPmsLwZcTe5mTFPuxooxoXWYYYOMgX42mAo/TlqQqBaZ
Ipyhhama3D6bz/2n1Et/4jD/pm3wyIN3LTkg8QISYrGhTmZgMgm97iFPm3646Zc/JMmUHccYAEGH
LytuUlX44n3mIoBklelzOcoP/SRlL5upx3EcSmV0SuT8VfkvCBBoRDaw4ibrnBYt9jTWa4bb9UeA
RnuOGgKf7JT9X+9Vpn9CgIuNVOWoXtABAH4wjs8x7wM5piPackPqrvAd3GcrDu2FBRDcUPducvRt
B3am44AVYDrRx/4QPjBl232FfKXCgEQQIG7N+KjTBN/1zxa/QLbrE0nUOTMYLTLgpi608R6M/esR
lh3LmhB+WNDn/KIZeMuI6uZmR1KwYUn45MFlGFt/vwP8Can/r1V8aRbDFgAGjF2nstjKoieB7HZI
gQvMWSXu9ItofaBqth2FQV64+oHxnx1bBd9xqgDVtQQ0KFPnc3x4e8zWGf7l/b+Wg4jran3k0y88
8Jh73y6kOoltgJKbjxj03XXGujebRjpho8717KIR0lh3Ad1/IcW+7CVPc/VvB5R7P8WP6OI7MRQD
CBRn6Q+LNOD0jsiMyzJZAWWW0w/KjARnYJvLZp8x5zHTcl52KEXuZ5aIOiD/iKqxf9F1H0GMofuX
LZ6t1Iry7I2jHSd5CgBdiEPfVj4Ow4W0b+xNRG0koxlt5D2MXO1UkIJUhGLukQ36Zn7OV2J42jPw
gALn3sDGxEazkRyffho21Bi1JjWg4+ccMVfeCSO/rOBrXwTr8YvEiC+0ptKCmf8ZylTF2IIXAoo0
2JvCrZ7UeByn8nPGryv2e3dvXIutmdry/62U3aKMTzyc7wUsg2tBppyzIzfWjAkhUMzY91Mq5urB
UhsCK7TpsP/UwRV1Ye/oSEYG6MpjQyi5NztyzaHPS87ID39zMasY3wmjT92GtX/PYRZfFdBthiAx
s7x2WEEe3kHOAZ2gGnuAgJ+NprAHCHNSRUEJ1fIkoq7xpHLTCMHj+bbiZH6MYpTh/CSjfuj3B56/
Es1JJc7j7wCzRpt9TBf8w1fuS8goWsonuS38zx1ydZ0zEKCtmeb2NyLlQg9LbHzu9KT8kBTXMWWO
yEplylgv+EmxQNPhJjBmy/peIgBy9IrRocUUaZFvKVY5hE3aNlU4QWCNzFmoJSgeK0ik5dnCv1HA
NkATCvVXpJcs3ohhXkmIK1hPhIg/2fxj0UL/IgiXHxot1y/Q39c7Xn8ARZLFIsRxE71I/TYKkQWj
rMuCWG04z5V+bFsn2WQ9yNCXkS+uNu51IKGmn29oHDdLoM5V+szs6aOaVieID0oUCiWuN6wgKk9v
h503rSo8Q0KcScYJhXFtXuvgCTvxo/q/C/5U+RFKZt/t6QtjyQ4OVPFa411Fmmobe9zS2MYwmoRX
11e5PmewcipFehQaF4Lk0F2REQhgBTKgvT3+JVSH9jLegdeevR113eGL54QdS9CpTvm4rjeultW6
7vEPjq5LpbPO+Y0ceo29INq0GzIxJEYjwWUs6Rbq+H3RTgUGXsneMIUeuxzQ99gS/6L5HZWbDW66
Sc82pmh/IYLJRj9poIhFzX3yLJI8rjfa6PMlVxP2JBl0lITLlZQa5Hp/N7xAg7WUP1lh/7WpompX
y1ByY+XnqSGnxLLN13vhSyOZGq2WOL7hvqyomHol90GW2yRF8lo3poolpYXhnLAQd6ef10Dxvhkf
d7EzJTsuissRjfnKc9G4I3kUh9xL9iWg8661H/AZBhd2ZQ0A3OiFtOOVt2EwhASbJihmL0r1D3Hn
U+Qtacc/LgGzhE4ZQmAVGix7u12U+YJUYp9qnlx8VEmHLteKErQm9TusmRdjdjOzmDbAuHpiohmf
Jb0XsvQtvdWKRq/3wBp/9XOuLnhu7IBQXasB62iAD7cJY3uuBqpnhDXcUC75ZYR3oBLBpG8kGnmx
Py3UQAo09EJHZnqC+mbxJ1rOtoD9M6tW1a+nimLTSrDBmtcVfKKtRFHLuOIHWSUd0fBNW2CRZF1U
224DxhhedJgK7uHaLkpW+ebCSgoihw2LwIf8nMkEVuzGoQlyBWmtZcCMMsv4OOpHPDuD1tG7RsGS
c8YxBLTu0rfO8svqO7CvA64k/p95R/8yk9wDmQfR3ALOjJcvZsbFOOwvQEqije+zaB4ulAwRvG8D
jYU/rsN27Kava0rZ+ZFS1I6WipM21arVwg7LABKtMYrP1IocqXHFKdqrAJHUW00EHwyx12jHk6WL
3E2waeO1p2h4LULyv5+y5G+kuWyaXUBBbrHUXRhI7Bn9OsJDyQFph83MT4wI7fV30lKkw6FhaDW2
b81Yunx9pn/zWWVQwm5547RNz2/9T7U4yiP5CVLz2y7s7u3unuYZiNRTdykbVGTpITWipWgekTbJ
bvYHXjTCDm0MYJG3S0JrajbCiMjAg4vt/tQNgtPn0TdMb/vvINiM+eM9MwinBFfcZ4YHZY73Wg6r
zwKFN35mkIDgJjWzBQB+cjyiJ9fG++elpIuIb65rbKKxMEae0EMj7uvJSUCMKKft+iCaDE1t2Smy
kZKrTYBiy3dCXBWxvPC+0oWlZVXPj1gl18b3lAoJoo0oi3NmcSkDB0JW5aTSO8LGRG5EVF+r59WW
HE4g2npEd+RrLUuWJ0txBhmi3Pd31ARwxMmzn1qHlz+2fHmXN5QOZQarQ0CXIZ3ocfM5dDpyeGko
/EKuHgxsbh7kXSGF0UKybyVeoi7hhJtqoFsjnsqr+DvjcNA1SAg9j/qjm4TWsQyXWQHR/VB8/Xfp
s1/PT8TTTppE/+bYvkZ1XnbzN0yvFi4/mMKzVCCGi/5U/hTL+pOlHFe29C9NWonjZGVMq2wt5iuh
Y5zvto5aWsLAUYeApAOcXsFuV7twhf2wbYLoMthgGjePoU6qjCkjtzqAOVO93GCbRaFQkwzaznjb
fcXfs48VkrlOaTRIkbRJXbIa+bkoNY9hh7l9wpFvmRq2JLL5CrTKTguqCaB6foInlB1pghayPxGu
mm9Il2wCtocRY/X5TzP+y2DqT7yJWN+d+2ZK7pLhT1hCZ9PlKcA45cTLxu7r3ZIp/ZhIyL8XiR4T
o1ah6P+1NYzYrE7cJg3jnmAQlcDFTqLnEPzSfNVWl7x9Uj9vxHAz45g3DDoyP3+VNrFfWXlRtQ9V
9U7mdU6yVuv8PqTQnKb6YCULOZni7Fy5lcJfyFtaQTEj0bDlTlyGyGi43eoGd+v0FMVlqE7JNAZH
Puepf4tMVbMjiLMvGal7aEY8BfTBuv9x0L9+lGOmwWlAy1fzKf4quwAzXIgK8WgLbCCZ7eZAeIiW
rGhmH8kcoVJxfRUbVaAEsO5FlXAqJwcbHmlyX9fmkaL2GDS40Apkz+9G4+8+uPoCV++ZkoBSbprn
vLKPKZW5j5yPaq1Y0WRz0NJ5VmR6ZkOtGDDxGE0sFpXukxgpYzvKl4J5KwLsufNd0uWLyeJqNMaE
45c7dnvNDfV7lU788GKBSZjOgwTZeIzqAI2dMmcIQSWsr4ABMLKovzV8YCDsrVnc9/I9kDs/Pr1l
BCiGHTzS2WtPGVxOyD98i0BpWcX6vHWvuQ1/4ULSrTBVSB/GWHWqp+WNfZiDgY7vu8upBK9XGOmS
2WgTrN8tDBiuMhLkEroL5JVvkaE0x/jutSjmaN6xh6OBNYoBkV0XMvcU/wu9pzTLm42jFrXrfnCP
W7AB/YrziqpgiZzOddEMHVbEneUMKa3XUFw1WJIzkdXlYHzub4RP4sPIq7Tmd7BNvW6Fv9Z6JjMj
CewcgQgN57gnoquC/JORnUFDCbCdWg9G1v3U78Szt/EkRyDdBBVZ/LyWybO4XH9GQqk62pYO2ASo
9qw79L2YaW8J0RjkVXN0/dTC8arNhFjR4meIdXPGj2JyemKD0wJ3r7vNdGwUSYQhgj7YSqKm/wwo
+ri77yIPUO0RuYxYZVvys4ILRvbi/9DJWTcVvJWOsNxSs9eeQjTE5AiivebPTMn9uIEgkxnu7vgW
o4JBhlMr7VI2Xyfr3RyI4yxIU+RQ2pcv6TDdUZhKmzoLeHJKiYoJZR8HJl/IEVqBNrH1ILXCpysI
YKN5sUBoHbxnpry4+8R1oODOvhwYWsiEZGNzrCJxTYWN7TaVixk1qVe3/TTrLR9oiZPdr0LtnQXB
SYpNTOA889Rhbts0Jztv8ahTL9AKxFEOAOqG5ACE1qaK43y9Ikx/76nMmdnyxa45Y67LQ510AxTh
xCjUC8A/TVdjG+3jW1LWeWmyz6XX/wk4B2awleJIhdudX44sXG3Q2R7muYWxiOJDetqDHOAMy8r2
nQ7MSDNc4teoO6YsCnnUsRSSThpywcvO0rBORJBxvjwR3HK+vrwnHLOnsnkDZwrExsmi6N/vFhe3
oJCiWIAQ/oGY9DrpOa61PpRUK5yWc5IsxNy1/0J74o0IS+F/a5PFgMyC9etj4UA8nW5t/XXQ2Pvc
4v194n+xSl62jpF8STlUWyxN8YC+FiqlGEwqxEXNcZY5YK/9nBJEfQkx73lbOSj18UP6QhB8sCI/
Oh7P9aisBortiPIDArRi4tf1hgLjvdTsTXaCayk3LZMbdKrkZeEnqRv9ZF3dOxCvTLWt2bS/3cs2
FFoGlOe8psZGMvE4I63gNv49cnQfj/dGBBTKv09mHLhOtAfsSSml+ymrDTaONK4CDcVEFxPSFooY
i5PP/nv3oVxxbJDUwLa/bsqsoBik699YdopjCHxWF03RdEdPAyoFc1h+/QtNaUCkW008aFUvZnLe
csa/O7nqy0HmfxlfmuDl7rujfQTY3RUrBpi7ZuNedE8ivZVZX1qEUpqd1URHH+RKzF26n1ktERRK
Jj+5SSeN0i6EZiPnOITrjtgBPynlW6ujqbJyBYDwBz1BhEIktQjc97nXmhadwRMq9EIHVHeLmeS7
JLqPGGqn3C7RNrBukSF3pb/nsR2fFsYEum5mZ0uOXJ/J4JaHiO91cbvWp1GM8Hr0NwBobRMMXisE
MMa7ajrAEWOvsNvqUJ3fR4iYrwM7Nwux8u3gu4oca/q7mIb2BJhEhen+QcuZf/fHiOI8tlSYufkH
P4F0f+jDhifEvl4u/QUE/m2wVrFCeuTJsS1tYoBjuswYqJCASR6i7Ut+GJHqVc3XZ69C1Te9thvj
jx0t7RfaPU6VqLVcbTgRCQkJ7TsdPzSkin7wHbZVyPJlCGlAAI+Tqx9IzEh8WMy1CQEQAMbyV5S5
Mu2b83U5PvZoSHe3LFzL6v4z6pnWIzZ2LTrxaDtTlvYA3A+0uoc7ZMURQRaoyD0YDGoOvD1kJJeT
NG2w8RQU+09Em7VzRxx3ZIHXxUKozhdW/NTQ41iDlqfYvxexQYAvqXx0ErNFj0OQFvuYg0jYj6/4
Lm2nenfPbZpHYuZIL0O8atJ4SPm1aZTgcHpvt9s2CTb/9zIWPtciTo1zp6Y6fxS/gBFmNR623oMS
vh8p+5fVD4zbj3vKI4zQjYSv8+nt3lHexrDRbwr/49wG/XAHdmqalztcC9CN9sy0npLikAPA1xJp
0Pw65oMG92lm1KcjNi0zgR1voS7XiPfdexlBplLRcQJkIdYP2WKwlOwaGpM9NXb6+l/bi8fabCCz
ibd1SMOs0LEPyhQCCCb0y77cCGAeCXRJD/sxWGbE9oLMounU1JhrWnFQhlr3qYSMba6PGyx1YoEU
uYK78mtxYu6AKTxoFbrBNkgc6tJNYE749CVDmb8msMTPBXSoBpiNgoSuDl5GmDFLQqQKeYzi8vOx
mDWvflTKhYxfBPmLVesujJsFi57AHfZTLPbFXQ2H1Ohzy3Ykz5OpvGigUMgn8Iz3veJvs1rmGnkP
kp5FK0qtz68t9kS/b2x1bcVpii6X9IUDUt1zx332l+fSOFCnwnLOdV8UWbXuNJEl3mLlvz1ptP+T
jmPZW7+pCA9yFzXflHBWd2Bo8tDlwxqYmFRCnSUMVgZqiBy/6V/mdPc8LSxIbu8koH7QnITS+URD
ZYIEaOWBHZJIP5Bs/8Pik4/Be/FtkgIDRAuARiS5k8XsRISKMXVvcafIFvPhhl/zL50vku5qwpXz
ObGrorr24KcplYXD7LoaMJl7t2dfrj4Cs/Cn8pVBPQkPWD+IkJwMqErbKDhEgPr4ILp9gRIs0Xiy
Tu5lj6oztMuzHrUD+O3Zw5Qri/ggFB0NA//7VySU0Kbe2f5e1pKY5HLB8smcYmRDeOtmfo4ItT5M
LVMcfyrk2Rw4+XBXLm0O9PUFEd20Kolp5AWEYniUx7CV5dRktEhsj8At9GrW/ARrciPiETNAs3ab
VplxlpZ6hdvR3eQ1zCDHsE9eu8sBIH1cRkSsZ1DtL/AeV4C+h/dWWLNuJ1tbAXI65oqPUYnqPAcN
GdgoCFTKf2M5d3OiaTRqwxHp6J0ig8QAY+zUopiPduyWNe/kwHpyEcw7v8JHiyOQcFXk4t4Q6Wiw
lXZ8kMldLa+uWXof3sIsIwqvuWWzLF43TR2K0qT64ZoVJtFcgw68oXynecxFqamhD6bGm9UbpmBh
Q/o9kv8RQHp4B2J6MVm05ycbFftFFAee7NGvgTiojA6jwiEZEWArmOsErVqhE0++yDLYA4IV4TRw
PnsAlcED20yF7kFWME8fldnyao8yWaG2FvUjLLzcgnn09jBaJ7yZqxniK4ZI4U/7yaWHwsrASoXC
sPeK2TFBT4EmbfDcuKexep7yV1NNyIFzkylvfmDo/N4eX43nwLmAfePGU6GnjkGBpHm2rfoSaso/
iM6WR2MM6qldl8XxdaBInIbAhdEu9Nx8LTfN5p6L9fJDx62G9FuesS448qMGC6Wk3Fg8UP9/zTry
ksBQs7LyU22kPtCDk8y0pn56qyVkN8mUoqZOFq/VT7+lzoTh67ADXkL+JRlEXHJ8Fzgox9V2926N
OTD8qjYT9ufMTSs5wktOWqGWfCuw5otBm8iCCxxTl3FagB6sQT7QhSn01cf2fc84ScLUAaVhXKbq
6er/yEt54qpCHGfQ+z8HWjqNIqT7OzQ9dsoiFDjiPC/j87PNpf2DZ+i4Ao+jfEFhgENHJOLnoTX2
EFa1kIHHvQXFmnj3d5WG4kizIKCiRbHs3kkhs3UsLVzK5tjfGsAxLj9jCfhMtKefSk+ALG9kWzwO
NVWqv4np2M0z+1sgMDoa4eFYC6YB4+WAKl9wlU3FaqgwhFOl6hG3AxC+tDK7yPYI0JWh+XkUiVaZ
1X3xmR4RfDE9ddtbdbk9+u/IQpy5/yFgj9am3kngC/frrBvXiCByai7RIORFCnHd/NcR5B43PEo5
eoBAIfFlqLlOYtCPm2sCW2/nrgqo/qPUuDTBZi11bzKdJjBDg9nC/tffsTRks7T1DbeR5H99Uu2P
7S0SzXobOLzhhyXYQtqQVXnpqsqN9UuIl7epKUT0xzgVReT/3YKPK4DAKyLdUOPirl47IK+rN1fq
H/Iuwv0ynNTq/P30UAhXKyL3Ud7LHtr/IHMUS5EGN71qC2u+Tib4UZOwLAoTClB6760h9TTQaH3N
ZhKTr/VvBmqwvjvn+bCpcou8RE9BSw0JUPCAUAAZpcCPWykU9eNuAW1haIMW3YJiNd3GJwSvhUvF
hyuR2dB1H4nPx96fsi/24kmhFKZc8nUSBGPC9M0jeL1+1Il1KyLQ3LVkTtDPJq0uzbdsMwaXNSqs
YVUigDx+JTadFgyCZOAp21AKrFGl+h9Q21xs56DP/+3sXjkPXF9/S8YjDs58+i42aR/NfCPlEIq4
hAIJSV0brVwyUi1TqdKjBV/XTN/RYnRwwijZs3mIaQtxdMRLtI+qhyHQOzwvpTGWZZlRAjbYce+2
WuMEZ1TrfaBHr61L5nUXuoDjIGa5134tQ4vloLJbSFPKaeY9veisQHc1IsfkZrrdoM4fCujhXym5
gBQPpxTcpT1nSy3Zy5UMD2UECAc5P78n3UwNJOhVsllIadFU0hASESSNvwB+peLQKwipaKQwGvn1
lj2Yc1s8nw0brl8fXoMQOWbGEWdx9tAQV0OFwy35WUcEnFgTvzzpC8bKElWcFJ+ew2Rg7F2UB3as
6jBdB/K0yKpmDVSAvR+FaXQQf7186j3qJMGto82s3CNrWHI4t9iPqeLaDfX54p0tt+xM5GpWyjWB
lBscCbZHXz7MI2/1juYzmtvfa8LXDJuOBcdJeayGvz6slSI15EaXaI1iswJI1gw+KPB/DPaHHlwD
Iq8AuBSIJlrD/LUaMn0rfiqrf3PQ1NtKpvVwZBEnHX1Fwwwrd6JveFaoXeLgTKC+De97+Yb+Rycn
plkNB1nfymQOnGIv8D+x/VTpGphx3uN6dzlBYpp1b7WynknyNGhb0pbhga5lmNWjsOg5kVYYBy6A
CewMd8I6RiD2f83QB5WaWTKILT/D2bHrfq8ep9HMKzZZaeUwD+uyX8iOsJ+GpbKOwBkmZuNTcl3b
jnQJ602+JxZlUQz9Uxhiv7hp9eHJp+caD1gWpOBkJADDXliBUkd0XaTBSGyauGWzuAkst9Zv7U4v
NFVokL/MpbJD6tIvo6QIgTMfKmuoNKgSQ+MvzImOz4Y9jVN/cWBgrwm6nvOjP4m3Cj1dg1LT/1YR
O9VOTxhAImSxOIdbofkaK+v9GDoJRVpQxLEPAC6bpOUgL3DPpOwJiolPGVuh6WFh+mFvKRvGqvlL
HkyyXoWz0uoMKcxx4Rah58awasFdQjPoI5NwMDa6N6CAO2PH2Q/cLeCyiOAWMWRlmsziIC182JaS
hZajPiX9xzDe+qSFNHpMFwc/wmeyfXusawhElrMqbW7Nqes9DDn5CxHgShfDBH9zs/AD0Bg8QZ/E
UHG99/wcPdM5FzK2fWEfk7Zkkb5lwKI0cWfFQL6AcktBUd70O5o6LoYdZW8OgW8B2W1R5FBHVEvo
dgWDZjxswZv9dqMBKIp2VfJXPNDe32SrVWa9EI9aGFa+XBBIWyiBxkcsdiJHcnqMAyfN0zyEmS6n
Ia6vpv/qPBSKoXaFPIyw+fiVCAnEhNQr/RePd07nqwRZWLPg73mbV9NW8kGGtPmISwQeTjZYxqbZ
0HWgq8lfpH9tpI9WK/GhJAPEJQfL8v6CNyOlZuTxd0vXMkJAH8YYxs0dgjXTVkuu7BdlqwZimyoi
3QBiuDf/gchZBehqJRIiqyQw7Hq8K+AezxISWGq9pVXZm+q87i3DDtvbSyTpxa1BRPi80YIlkoxx
Zo0t12i76wAoOXD48XK0HIogfq8p9HP0KLWaSVu2zCmmEKo57lD/RCNP0+9n/NNV/XlGSARfldnQ
MchNw0iTpIuCy22M2ZzmCXOBLiCdVmnOP1P7ehWViGhDukT1tlKwqSXN0+GHxibV9fJ8ba2Qlxa+
DdGTQ/cXeE9NRi1AUh6yT7HXdmze7Uanlgihw68cVOYyjVd/i4dRULZBKWmgkqwWWjXKxwyYkLmo
o77M6Rbu39b2gMixOITTKWK7H28aEyK8aFg8PyszHdy/orykCApIEUNcDNyAgj1m+2pE4kCL+3uw
C6Q5MM2jc9LQYMynhJ+vaUuu9tmzgWqaI0aF5Q5EIQ2jzD7Ei1kXJgqSfBjPaXAKIZD/+Xi8Nv0y
j9qHxgBeve49Q+9GI+Jc1mLSYEg2xs7ssDMfMrKsSHP4DtDubHxBiKkByoNJRqTF5MzhuBZDKOmH
BmvGnJwNaAxWelWswog7/stAerug3Dy6pHKP9lZAspCBQUY9hs7bvb93CBuAJGtbzragSaKxCkhS
CJw5wmEL2cpD5nJeAL9H9ccuYn782TSPn8MA3XsL/JINncDTmmXVSuJrzkLvpy9+Q/2dkqfCepoO
tJlwQtv+mte0X8w8FhjJP9LXaxowOAsOOp39ethavo2N7tvztiTWjbh6J3eGQVtM/pbBe0ETXKnD
jWxBOCvR8CNAbU9zw7t3U/Az5PGxiKmKBx45nebhmAMIPzOaKHM5a7yop2+GjS3JsFOqnKvs9Ola
U08/QaaGvC8hUbWK5ReFk0t/eCuJ8jofRYalWqLpmZ12HvyCeQ6ylFf1dk9RDrDLhYqAeaCYD4mD
TxVdX8yW87lM3/fn03aH4FtIHEsUe7VNc7XfcANXn0RnsBZ3CJDm1vIq6ycwwLBath+mki+Gprau
33nl7HGSkTg4ErMjj0geOU8kYHJphtuQx40t6I+MsYaS6mqkm/GKoDUuJOeXYgLt5XeR+SVhXgaq
pMy5qfP4K84OrYiKZZJrWdVOb+A9dkX0tCyv1VrzqmeyWiE3VSBbCHOBnELfLpbsRbYUSbgcuemM
k9XIa1FucHeg769IjCMyk8B75QIDI+TA6ajb93zKwxWmFOr0wie/5rLOBjDMRfs8r9b0ljPwjK4I
52yfc1lrVAfFqmJVPUUTKHShW/IVldedI7qn9Dvuo4mWL3vvVaBFfzgSBOCbjthecCvIcm1Kom72
i1+XjYfwepB4viMozmqk5Hdvq8i+72PhuxpBFi+iOUkJwGnzfd9VQqC7yF68sOppXcDUm1/FbuZl
YKCj9F3+6dtQbfXsSlBMBBDz3evIlPzjxbwhjaTivzDeWOdkEX9dS9dMrqhTNHFVvNVjys0hLMSK
uPN9OzqCQHxJz326fQaVE+RWu+nY5OKuxRvQkQF+hT24mP9y6zema8Mr849zICx1Rc5S+1Nc0Zxx
yQyznhoJQLAgJc4I2rcl8POH6pRg99W/oYlLPMQ0T0Je4lJs+i1C/7hXoJegqsIXwjTh8uZVYSz6
AXTuyg6zBWzw5SZBACZnlKhrN2LK0pdy/x06U44oHYqo5MhlLDYVZVU6SMjCk+TZ3ytiJP0c6z6W
1wgYALa1XLUSV5OezyIOXU1Cf6qrtofwR5COJydj7AASnwsVLz6CrwiboZkw5NyacYhDhKJosrNS
Miwh984zZ/0SjC/27OrjrQBlPcsc4dHx465a3jbenNLHkhKGoL7BdibjSckETsfr6hIN6d6GYcli
NiIoPis8CSXMu47BtzxII6OwX6enZqAneGjsXWFkk8k+As7ujWN/g1k+PpO9aAc44ojK0pMR2Zdq
neIvSsKRcmV577cnFV7UZ5uA2KDlJxCeM5gvWaSmPApVzwC3+mHRfQB5cXtN9ZUs2LOq8JzZzJWD
7tnDann/l8kdV/w4vDOqLxMqTRbBxMJHYXZfZ7hhYr1P4QLyglaxtvJI3C0vG7lx6IpVdkGGThO/
Cvhg+yij7nORxG1agGQw7StrE4faB9ik+EJOJlBZsEWz3pu9WiLeryZp3zMdcphD9/KL56Mz2DaZ
+emdcgfIuDhakkFo2Rkl48XqeBab/pKZ7M0zH9hb4Hxjt6wHzlro0rj7SiXwG7h818QoffqTrgIf
6gpJeGwqz3XZlDD/koymm/P6hJBM4s/NKiL48bhF4z0h293qkZdNCtivuU57r6825S2TGWyVRyFO
zsKjOE0F93OdmhzyCHi8QHOPsjWq5FJ2UytKSoVsxqqin/guLDgbuOGqpMcMt1rFrmrHq5aHuGI8
Tm+FnjzDhXo53Wo8aB005WmyBIJocF+KAwbBM0542+M4tTKIOW2z1wZFDeRGE4dA/DTSlWgq5IV6
FTzq0rf2G1GhiZiB0NTRcGYj0XH/gPFSH1dokZIfjpviD4VEX1ETU5Pgd6wDkDrNMHSbVnE9cijg
SfMO0NHTvqOzn9sERj64OyQOux6Z2JuJmIMc9zpFeIj/+pWgaxu7K2S3su4xevbh40gta8d6he1g
rtRDVNS7pFTocHC+3b0wwTX+eEspeKNo11Pm04WJG7SDD/A82Wk0FBM93d3y38oxJQ74eoB3akVQ
WsGW8y7skEqq2810wgemkg/+l6DuEd9yeiA0nts06pY4SD17de/nEhJcS0Dws6IFt7dn9ccH0CrM
EgBI1zY8ZQ3hovuSCPi0HYHYBbKm8JSXX4aOK99nZj2/+aeLVBTnw3hZR1B0yXDxsS82X6CT+8jp
81rEYwM/pLud9Q9SEpTuLxUijjpVdhI2g461PAZzFqEMAP4UaXVCtDLm/YwOWP+5AuksMg8KUzXM
Rs1h/M/sHoDz996O9en3I2yDyy9tMFxWRnC/VPFqnFKm3T4UFNNpS/wHYxucrezubaMhSiN7J9JD
3OxPjs9aTfgVaWZ3yCOmNaZKNb5uJPKez/ArQN6AR5AG3l5XH+63tnyauijNZCu3ilVKiSrsT278
AAoR3HQzaayV3MO8L0P3+dPXGN6AeEWYJkMO+jHoq3W5zsLexbUDDX/Ghlage0oyUmUgyXzzjEXo
hGJXtS0fpKzQC0WRFYSnIVPLDxeY4VVaf88VJMTS1A7BhxFa/9bAWJmVgD1+DEEXlUeXXgz+3kZb
jLhI9TL/1kQbxoBea0M6bgY/2pQc+8pfRKr+M7sVcwBKivbP4Y8AC1tbkW4ZpHP/sH2yH9ToUTWG
OdDuFr8q4LUkbQkjfnisVnbSQfaPq013Y5Xo1exAnMxrOBs7PpusAusATqbqw6eYHmvk6qXjxk2A
TCfAM1Hx09l/PU0KhGWFBqAFirs2r16eYOVDviUklZ3azbXDAeeCsawo/J9qy2XPdt8Zh1cwflC9
F5BmMD3SRMt1isKKzP8BzECbylK3k6cx9Eg3ZhZnmmNARz/kZweZ+1APshjKrhbgft1v6TW7aOEF
jz4MbSQjKmoFB18//UVsgw47uwyGAi9CrTkRQqlXoj2SXmsrv2pCIkvyn9rz8Twqu+wR2aDC1C7h
VRENB7f1M6K4etlvA7A/7NbVdgqsQpI5Q9pDokLYnfw8r0PIQx75K01mDU51VsHGZmKhdciCthfJ
InwIEEmzLm5N4aSAIiMN89LIPAvRTA/yN3wajgTFAHztFBhx+ACNasL3/Y/C8pYJNhfbiu3PpeE6
wY9QCRPNLOwM9wq9u+EkwxdeFA7J6tkrXEng4fgs3o+OztetvIfIGH8EoJv3/Q5I5CjsMregT34G
3QGKPuvEgtR6t/Tsi2J3rl1rBVYhneIuJYBmcCZeTNEtUGM6m8cGP1SX0lyB9YTuDUMlewlJKIeQ
9fWSi9CmQjZWRWfPkhYI6qchhBUhkg3FLP6xykQW8dQfW9GxTS4UpSkhDOzS6oAC++RggoHJTCIe
/HSwh1EVGmN1VI5V7HN7jnm93gxAwzYT5o1oJXYE7gHXegsdkKNsIgNTVJcOoMSS3GGlSezjke8i
7kOCzpz/KwrwZY4jFjGDMLXBikrORV27RE+ISS1Fbnhi21BNie4ui0uE3ZwxY72gnrUmGizumwN+
/qRZwVB69iwZRPaN01tUDop8MfZPL/IarCr1EXWeJJL71SUFyuZUNdkPyqWnV9FQQKjJk87Abz5r
IeB0P0+Y/K51fBdbg6c5x8O9wimZWeFg7YphQg2zPNeDF+Fqz6soq72WsCb1r/NBRnOL3CXMnjs/
bHD87LGnRzFmUsiNatWh1Da6T7mNmrYpuFVyBLWb6bbIjFoqma5ilMzbGZ8sJKGQgG6wrm7PhojV
1McG0zmOBPo2v7gqJorJjca1+fuuZAC1sH4AqAh0/Lw5Lc+5vRTWoJYCmvU7oAsPQLT1eNYOr1rx
xQzgoTgSdS5IdEKKpsIpMdjPYkMdbTJkZMnDnn0nSM8JCvx50WTIoeDPjrzv9ZloGschjaVnZTpn
yVjjqZK15upexRbMHsaxiS8uIwFTQ2IfUlDgK2ykdcBzBjqBtJ8JS/Hqf909o0T5aJiVLkFoxT9v
XDcneP08nRvkM6WN6sW2c6vQjMnGFAN+LuPSCUIfMhpiVLCCem+F982qV+SGHLd+eA3D3JGa2EFv
xbejDbxYa71HMLpy1SvfPow2EtPUx40sxO7nHWTat/EUw05iPEago3IxpmSSVrmpqOFaTR5P+Oin
h6Ho3bBC0wmwZXfeFhJpAoqvYJirG3ePNkkfqqpDs6NvvIOuyI8BaHQBYPczxeSImi6z4W5QX3Z9
i5CL3TE4XkcBobX/4gAeaVFHw1w+yriHL8iK9eWkOgyUck1dojSA077er0eEe9d+RP29mEos+viM
Iz9I9mUbpF/ajbpclmJScQWwavBc2WB0kMYQ70yOHWfUXrKaq3BJfiwCk/oWOvDtGikznuwI0lsL
s4S6HVZ/krChzIarJsuCLZYT0TtwUmKSgYGzWn7HtRZ3Lmti0WmIRGGrpnOYPc7OsK8jta/rORd4
oUhTeGmKz5fi/RrAQkGCUjPIusFaRTz9Hkr3gVbay+EXqGwiZoP4fAv1jRUIN9R27tUgCJOh8Qk7
F4//OXZeGENjP6GvHIYo/HtEKfHB1JQGf7yYZ2JrOF7EPfOanJiL7pBge/RZ5fL5Y7215MvjOHRP
SeN4sAtcLQfzDANhIM84RWLTkcGlM0qScWBaiXp8dCY8xNReXcie03DTsbTAmCmFTI92YejLTprz
DvpY2rLvorSismz15kFOySRwnNSIGQbPmbymWnhtA+o4aSeUpNG5U5GyoAAcHQm/sNHgDl/JTCCf
ebpiodRYKmZ2322XtOkqjBpBfITt5SigrCGccK0P/fVzv1wSPbx6FDRD0O98MJ8zxSptugWgKmbd
mZj3C1zazLQHGWNZYQ3IJcEY5KhyibLQjV2pR35D5t3xxFgdntAIf17VWUniEgo8CthZTVgictfW
jP1DHmr4Ag27EMRO04ZC4sN4u/UKVfqgg//3szkzHIdREvU2KopICd53Ssvg1mC0HHiRfq5p1p+5
FwwfTewGjJb3/JLQR3Ne83Duc4DbJP/tkUK5vNwaf5TeJXbz6CT3274NdPsFvZT51dniTYdiY+PW
wQfoQYwrPcqg4wnCcaxpC2uk+DVRkdBodI0dTdKrmnueAaXb5vOvbXgY2X4nHXAiR340g7lrcd1u
S/kqr1TK6jQNskLO/0jZHn2fE1sCs7ln+68HENLCpPdwnbPB8q7hfZHgZ7fE50X33WPHJ7mvEJt0
hklmT0GTMYDmY/i+qy4CvOmzLQRdnFheGE6kcMkvwGR60Fw6gG/aQ3zFYNqlH4q2gLmV05qxLbET
RPKpGFmGYa/G5DH25fpSU7xsxoCkFs2W/glPuKBYTiUOOyyY6MlRdIrgSp/yrhx301x3maB+kVZl
jrZDohgV2LfrIOFPPX5NWPMylXOOP+S3WczWe/FkIL80gTrZyjQEyh5vNM6dnUJW2HaYADV1nman
x7OxXzeSWB1O6dGWOxx4u82gM4zJJGi63pkPvtekSyFGoi1JmQbtniU69hKr/xbVb7hx5VTxz6ae
WO3Uue/0XC1+9kPvgLLfsA8yEbgN/pm9QLkUPXwgjPVQjRC8dMxprCmjoVBbQcR24JUD1PjmjGqX
Mo/7tSvwGOzD4P74UMfrZzG1nICHkoSi7PIP60HQ5pjq9D10C2FTtMF0GeuuM5kDgI8U59l/XY46
M/TZm5vs4DpTCp2w7UFyqhagUOjLSMh4uAXdBApFGVshx+phKR1eDtP4nslr3RfUIRjs5RLLGroe
smqSnJVezVuWRxiiLESvc72ZAQfo3i4wyI/kBioTTmto/yKDIyXDdAhUU7ReygJyY56reU28VurK
FkGMBRoQ3NUVB4PKDUq74uwhflsdN0+BU1gaQy5jaOmJCMGa5cz7OKOOwjdmT4jXl6TG50FdO6J/
jWFqOl4hEPY8Ae0DKe6hoQescZZQVEx2mNwC0p9ZsfbSfFcIP0W/bHBEspDrp3ro/tdfGFOS2WCH
eqyXme27yXwmeQuotq5WEF6bm2jp4b8rJkoRtTzidC24u5Ei3tcKsFHUYOJb5kr0h6tKP8wCfD1Y
KLpBcZMFE6Ugj8f8/BoVJpOfyLdwqQXOkluo0hwEfBWrDeKwauM/bALhH7rBwJPPwQCo+lhBMw2v
IbtIg2lENY2lUgrUSxqHxVKQOzHmnqimT504OjxvbnM85+OA+r4vys8OMaouvsPgryLIX6PvttiR
dFQ4XHa54VGG/YZyGbFeXQ9gbGZRHn1X5FAGezBV9Diw3fthH+prTR4m+Xcg44D0i3bpJl73p2IS
UdNq88e53KneutjPuN4Y5hvD4ApWUU+zElf9PSgdcoOHyQD9t0OMpuMGFhhLU78hxu8y+0JBOYtA
3NjU4NRv+4Kuruw5Qw1GxtHo+V7X5efasiH1gbdp3q/ddcP0qiTPCpk0DQ3hzWLLWCNhrMw9Gh3m
LW/Gnc1DqC2gGp4v4TXbnO1TC9DPBBELKnE+uTD2WgQ9Ui9EpQH3UZ4THvvFJctRU0ikm7AKTHgp
W2n1ue1nsXs0i7uE4sEhdB6YEL7FPA9EGxOYHMM1ftxv6I0bsrBMxm4IHwNo9NAQ8LePYBaPGYW/
edIeLAOZWLCZjv6EGgwPzLf5Rx5LFD6Alug6H4utpvnVfhGCKKYEWA1PhHbcwSQ/Rox3lf1mzYwk
7NG3bk6MNSvAQPHiUEj01iJDlW/LxO1BOw2GnxAnsyrF+mNfA/YcIR1G5DoiEip3Z5BCXGqIU6zz
EC8qtnbEsRO4XBDhSuNaJfJa5os7oMzs5USOXJcfCOCBcK2ojrHNhrLdaKKdw0DaDS9kfR1eODEq
c1E3A3WybhZREohV5MiWSYY+mwsRP3ZK+CfHvfAiL64diO/Rm0k27Wneg+IIDjpTdNhxyR4sY++n
8KS1V63Fmg0d8HpLqRiAhOB1F/LNyjyXndmZr6pilcBlkomrQR2DYNQpVm8irsB9mcgnwKwkBhVA
Ovs5YWTFbKyAsUpAiq5u+sOBFVdJZ6xDAyefLAgtHC1uCAX4Sf2a+NKVmLNZpS0vVmYMEsJVHvvc
WYyekQQnbCNhhKZBDlKEEWIKVN+/WDLijOmHMy3INyu1oAcVSqJOfGMUHpGQBW+1fhbRN5NJ3aek
i1y3UpWCWyAYHZwZZ7z/90FdgNKZCu+I+yECv34Bkez1P5pYkyovtQ18x6Ez7XBKugYfpBXAb2r0
pLeZnJHF0v4b3CzlC2Ru2RnFNeytsVs2fvyQiZL8F/w6Z8oA3DS2E6CkILplc5L7b8iPHdj8gc0U
ThZE5lsdCZOwZW8o7lEs2qois9BEzFJZ8WjVhSAAOq2Zxg47OTRHT9AJtbWHb4jMstzqUxMxNqIk
uJ8IBT7y42RRz5d5DoFPIGZgPxpRv9aOkOioW+L6EOy9i/2KOJ3EMW3mM9Zq2UgPXd/ua1cF4rkz
Cola3sQ6V5PHAEd58OTm2YnwzVs9MWaYCoYXKqidSuR8njP48SZ0XXE5N8Z1ATHzyOTov8SkHowW
Lt10d7FLkG70t4K9syBA3/vWaCchcZbgmvn6uejhaDME4X8XWeUXgSqJ3n9xJch1Ukm8Rc6Ule0R
AgOQyY3HnFISQgNir8cKWoZ9kCULdXJYVefKCPUXNFfJSuCBGbw7GF/jJsTJO0nk2g4iB/Yzr5pu
oMW8c/OjNtgrhPiTstHP6g+SUkw8u8+GFjXLJG0LlFa19nqWVwrohOj6Idfv3O4pEWygvBveu/M4
IbEYBSYxueuegpPEjdjEkczCR6FM7CKuWYrRC3X6iO6VGB1IZQDDJbYqIFP2G1RE1jqzKkWzTkAP
SDbNiLaGxszDSS53gTQScVL95nD7b6SejqdPblROCcY8P2Ve6HUnmYElubuL//f419Z1qR2cXKIk
uBBR0oCQEbYWcaxDKMee76XA0TnZPM1zuapVyHNLUZxnYsbKDYt5A4zyFcjPwXCfdHIi7TepsWai
1tO1o8wgvEEntXqcTCsS2lnnitDhz8ACOWzD8q76BvXdx8jzx7qCiDvexWI9C00gsWvOgev+t1Z7
gKunB3qS15qrCCbw1DQxQV5VYfOLgEl4i/EYRENcvRV++540h815kW6rQ3/fpPfyQS5rX1QgOY0z
YulnXtwZunpMiftAYSRD/pjrTsTBS4jHUEHBx1DaNKMc/5HqAfDBeRpYEt3WxZ7/wQ3lTh4uSSvQ
vZo/K/C1RFqVS8+dJ/tzfzw2UEGyrJTZ/S+WZTBrztLNf9wTwuf9lrLKK8tHj2qUl2PNH7xyB41h
Ew6YJ1y/aRFlY0xFyrMivN8rLjB4RqWkQyLAfQK1/zpzrScdwfx9ttQIjW1sjoZw6eEfxF7SEljk
uX+LJZfmdzOWnJbW9lnzAIMKvMuUl7HtbARvAMD8Z0qbaMEk/RQJlCxB2BS6yleOy4gta2tBixCI
p1UiGGmPBi+12jrWO8FAh3efubhnYGTuTM88ppzHSB3TId9SQxMhom/f2V19mO9Oqyrrxq3mVhV0
ycJQ7jVk3OoGJG/2y3kb/TiXAO27p/jyQlgt6AA5z3hw2mwwpgbm/iHAd11+KvzleChJkTyli53h
P86SZ4jsLXBSncRLvJIEk80YGFLGg/UBUCJGATVESuocSGNVm9Hkwwt4Piwy/m+zhxQkJ/3sO4oZ
Ea3AoqgWSjJ5wVDwKXS7EDFwprcUMBJbSJMyXmuZp2V5u+LXIGksTEvFjSp/VImEQV7+Sxd9Lsqx
FotFg6qhFtKUMCAHnj+XJj19D2FqdW3ePxox9uiMvL8uOh0CFuJrfv/icC30AOc99FK/3TICBuj7
38N/sfNOVKSbv3dmRWG+K8FRiYEVxRe6qIbW1NdCyGcQcP6m2+rVcLPJVXG9vMuyukR+mb7Bb7Hx
BDXgeFcRH7xIDq3MMZJ63fWGOuzfwxjpn0ExM5ENYqYZpR59FCuh0yWp87/YtLXUcD1phYnh4J1K
cHIpPlAl/JGoJq9i4v5BpbCejBCWhBjS7LBpT1f3TQfbT2iDCTj5tJoWuAhil1rJAX+SUPyNqoTR
8evxwqrpNhH05bYw/SiC3/qPgA55epStSVjzpSpfPtc8JujMicpkxOQz4qK/eNFKOOsiyycKC7oi
TYZFnwfFznypWye5vBd9WZoI/9ngpnkJPiN/A8QIDeFlthyThc2b0jZZqyHx29EJah1wMoRBkKlN
rU2C5lo2+wNJSqGecsJ+b85eIgJ2RCTasPkeZiOEivGkrmBdIa7a2g88UMtvnt8YXPKaAjePkuCy
V3SKJRtTsJFRLI5NnFp98N8NH0LOXTUi7Gc2uSvjiOMMnmiT54YIM2uJeNd41QlgvsuiZmBTD+OG
wOpLmlN5Kbr66+WbN6VtAdfU562+pRRUNZNRJ1SnUzugnjBuil/wZrqmVdD6kGgHFT6VnF4bL/jT
hEZPq3jlmn+0lIdKLj6QcZ8AEgwH4+CEE3YOeDTravjJ8uVAl9gll87Zr8pSm+Fi3ZohnQ+CJH4X
S+PBYoReNdPfkR/JRidfnYr5zZWfmjPfuJr+lEksd0VFW8GT3H9AXa9SBY5cN+rzyodygeMpy7YQ
r1EczyG+MbgJlH1e2glmUKarH17jRTqDkJFQrIt3vB12yw3EUSY6JLC1cfm8caaipsq2jhYd1uK9
VPwWLTLalnJCS99lS1Mjo1MAtldMAwUdmLPEoZFg1hdXFEzWoJZcFjFNw1jXKfsz/nss2khHEr7A
cTxw0sjDnn0U5eNSV3K8s5E4xGC1P/4mlPt0P1Yu2LIq20n/5os/etDymwDpIqzHb4tgV0cxuvX5
jWOwMzytn/AfKKJjPpvVFO/rCtSOT7BeGD4tDXNmRbk5cuVY9RgWoe3rCGTGWv7ntXxwWh2lAJmD
zXB9Xx0Kzf5BLv+rvmcyiiYwtd7FRQWVjwzF9ZE6+Q/o+xOPis3BowOirQwQbEIVT9tNf+KPWVHp
BdolSG9uk71w6+7B7DHFi9Dva+yRGOfsi+1kUsPPXYk6+cXJA8hrM3rDD1DigexqRkaCSCCmzbtY
PZ7uwSdmc2BX3TBM/scLsj33ZkhGePwcIYFuj8aosKi8v1uK58TvsNOtUsQnEbrYnyFCPo94r16H
0wZ6NFSvK0rwMkyS/FaOHTO1G+oK1ZugpOclBZf/CdZyB00pzlBFp3SHQtjlBre9SmjzeVXSTBR+
ybeYHUoB6W+wxJxN6ohwqq7KfxHNLsm2bWFIvW63GtXhfFeWzxAlJkafnTFVGI+6P1YO9CrJLxKP
QnrAOzbharQknDtGMnZb2ywvXoEuQqBw54oXdFkaoE9Dg9Ak9dXAdHAROiqrmYZBOKWe88ye9VZA
VpeM9J7l91MjxC3Bz8Q9DAfTHN4HIDaDcQJC9dmxmwrr9VzVgV6QGElR3MN9Klx3x0IXCTx9a/qh
SkxJcCoDTvmY/X6rL2phWPNOeNvYQU/KutAwZBeg6jgOv99XQGHY2sEf9omFJS84sZUfQOQ9sbvg
BDSY8eloJbyoA4bOUhdXBF4Kop3iaCuzqOHGBoc72iO7NWdel264YEjsuZDBsGi5li83tB7SPF7j
3gjCncyY5I+dSAeSNlbfDP3rXKbE9X0PVtlkj1Qnx0tUYJN9cazFEZmNXlGtkVFnqNuCO6KJOuuU
uifgF6I3vaoeD56+eH58p7rKXoN2sa7LvEpJ6Zklv8Wx6Cyf5QA5bLPJqdzfSaimhyyp7McB+54l
sXiuZH+CcCx8MGXwHK6ApzMvIKgHPEFAW83SdN7iPQhBSaEaUyt4HDUt9yADlElfkabTh5VdDO6O
OQUh8Ljd/hOeUwQsJjN7VXa3/a//g5jUYl8e2WSn2Mjj5mox+p1IHbegq3iwssy4uH3Fy3Q97OB2
jW9OqN2OjNq+E0PoGVantTwR40DTFZCRzxaduviWWHvwhbVHGHo5aR13Io0P0T1B61rF1TIPMo/Y
iZvZRqsW2dpqfUftlhgO0PvSEmidLAOBQxJiq8qj+6B++Mr12dGIL+3DtznQXT1jym0vAkU+B5Kn
CPAjrmd7l4a0fWVI3VXGfmYYorcDIgsqvCTg9whWjsx3z2CYGTqHhLUsZTMH+0bwrwhXj9LUyN/m
meGALDJnhUT0I+nO8sm3hQ5xZgSH+xLtYx5cZloieK8Cqe49e6S4Yffn/2Pg3UvhTcx8MujmM4Rj
kjeqD3FSKL2127IHIZ0XGLWXtZKOICfXvLSOunRn2NOmFs0byHFaK5P1buq+lsbaoJORrMGggtq2
AXjMHbjplUsNj8Of08+kXvxyLF0ucrCvwc92CQ50V/DEXl4VyLTKLXj1Pys8nHMnO6q3he6DRtdU
/MvGtGvj907JS48WvVwSNDITuWDGWgSRAT6GMUUIEHUdHHMNE4vTl9hcOyasqHJoHABtuhLv5AjY
iptEqTmHxA1YTLF56Yi1OdowuSF1NjQoqFYIQc2mx1QbfswMOho4VumbN4WPHlyypedW2OPMGYGc
CSIXHN9KLiRriBfSbWLM9ZiLlMF3q2DDw4Sc6hM1dhIqaXVruVf0jj3LwRAsFcDWYclnwHeYoYDD
KKD5oQ+XRHNSgjMJHSdSftch+MPfxiXZGxIJ0X5c6I2ttxdVjaBf7vJHXfkk6yKGXwh/7VGG2gbr
wEV2CyyUszdy2GaYTfyd3TxqyvIsNV/EilHhj++Hv0rXQY40ZLkbWUEqKtrfhXuBGRJdh1AqHyqK
fCLRs+pxcr+HcYNhlmagFBHw2knbHr63z2NGwNBvdrsl6H9DW8YhijKU8dqIBBJoJU1UZ1I19qJJ
rDJ40E8AxzLfNA3YWGCb/IuMcULQLbYg2KdGuw9MdYtEub28LJBX2s8LACsBbMhSGR6sN6YYCowx
I0ZtzdI6vBsCB+mnnsSMSYxlpWO4Pyzh+07i29fXhXgsB5v42naiUADQ0ci15z9Tvp+yuZX3R9vK
3ecFaf33HE1BjNT9QEr3jvbCRlInP33uSJ43WpIJKBGjPzAh4m8iGpzRxildkUf2OxFT5wBaQ+d+
5Dg7QdTsdGx9ZDPmUhmeleBEdCdL66hd0lowT/vGOJJE+Twkam+WGCbjx4bzL9wHeJsAndDcOcbs
7kUL+SuTDLCiyHB4HxtLe0LCi8pxV6rWydBkdJFE4r3yF0BSVgoeE0ViAJkqBlFKNaCARrVc8toZ
JG9LfpLNpIKG8eKeqhWsVqbkNoqKVVoAou81cgWGIHkrZh9hSWhU0sgh76vH8XDDe+oExRBB7d76
WUd/sg3qTyA09EyINRiYHKuMIwn4z75BE5KZEJ1+2UKtEwSQ3PxXInEdlanN21ImVgl/G5WUwusS
cg5dVVVyLYkIlbaeLfnWYfqSe2BsVn/fnF4b+iub2dEQ/eMbiv5syJBLIetS6dopE6C3KqQh/l5u
P1Pzh0jiA62ZuYoPuWWwlqF3TKgbj249MjjuWRBijFoo0Xl0zw1P1h1/1CKnaQOMygN2nIFNHXLe
XFPR5u9gKZXtUFoD1sI3h1I9DC7x9yQ94ZRBO9zYJijtUbHOciVi+BhOPDaIAJU3wK02sHT9J++E
8rizYUwVSgTVyFyQzXVPJ9Z7MZXkcPBHH/AVKZduY9SmbUHI7WrxOYatSWGd4ViNB4bg/p3xKXj7
M60QsYjHACCHHis+IaK5YE9Z/+bB0ETYlZbx8cNldvMsNbPyggxozDIFstLNs+ET/+mqyBWFEMgZ
j/ZLVfEKqYkqzBP+fJbzxeSAfpbZfWXJdyloeOormhkdC0jNMh7Kf85uXjOIO2UH8aqQ4+GD0y+h
x3MYNh+3NsaWc9XlWRwUJpOP2D0pFlh4yj3ux/14axOhIbcRBS5QOmDeiAjeXqjz+ZV0fAjqCH/4
6ZVM2Fk3KRs+IwDAViyn+M+7zjNb0FoE2kOa2RXGE7SQzXJI2Tlp6cGq8cFK3ku005Evy+RA2O0y
9GTFDnAtck1umVRpPrAmfp1AtasaQHsdE+vW9GzNwohZ9+tJouvODFTBLanDjUQI/OpxleVDLII+
Fi0BiDwSDlj3/DV+YuivjT+ozMjHJVRD79vrWZt1noJ2bJU8yzyBqXGy5tutQJFw+tGRi7xTBSCZ
d265iuUEJ3ZbU0iZQnnrOiwd39Tmu4b24LFOcP4FqnyTnfz5vkuRoz+x61XSxliK/a7K3eTsI+XS
CTgfjObWV4LHTzj0Q0Umn+pZBVMogIGxed8URdojM763DoEEtTIhm0c9hE150Lg2JIQcU2Jsxkf0
k9tnKp/Acm3e93Olze8/7XAsoav/ICWxzISpmA8aXEr6gs7pHW8lE1AOvAcLTGE216G0plhtObDp
DnANpNnBwIg747RkiSG/LQWJcLIN+oklQPBqnRxM4stbygnfkRw4yHkt1DbiQOha9VapZB6Sb3JK
fr8pYs54Flq4qmNGGCMw2jtqgQgtqfpEqDl6y4wnrMYwTeAeBqNfeJqn0rK6IJI92DAQDzWr8eiI
rBNck4dkM6AaRNJzA3c055VTV7dPk36GSNhIcRGKsjYxVVusWnri8m8b2OY5B0u1O3OD9tppWoCJ
gKywdNwX4x02nI74q14kwt4fI1uMsbXmS9db2lcvkuoYZarv3BBeOE2ojW16d5YQzyj6bqlS6FvD
BGbznepELV98JW3GbrO7kT05JTWoh8NceKk818YA0FPfnhUBNKR20XnIyjyNtNsQMdKGFjrV14aN
Mbg9/y9RDN8U+rQYwDogUC/s10+A0Kbiz5tyVDfqO0LdC5ywTwwFoq1xQ2sW5+tkq0nlBGBsfiGp
p2/0PnmWA2zD5NlBmg2WnHDoXPjsthltRuxmicCV+ueW9dnth0A8kzeLNQGbGgmifoeeAvzimJ4d
UoEWDLUHdMxl3K2o0KxNOf0PZImlEEvZsNMGwx3yO4EJd/E+1cFlYJB52GJcKYbITlECTeopMhom
+61sla9Ttq83+hpjyfiZWHBAvTp1+kffAKJnQmk5/1olxgzyt4iwPbJnYW2GC+Uldlj/vWiLqMS/
3Bv23HTqP6+Bz/BXxtl38h5aK2DFjkBSngx/OoYNG5/PjMR+5Lu2ZI7eUkyrs8IY/YLpWotiv2Wk
dadBNPsulkK+/PnAwx9WQ2GVpZpBAI3TOlTR/tqscccxa4UomQgbRAtXB6JcYlFvQVkHJhAEY7OK
MZqppooXi+toES5AsBQUY3D5gh19U9uoycWDfxJQW5d7Hp3xhTzKUElcDcIkvnU41ouveYTiYMu8
D2hkY8GbnCDVN2l949O5aV/Kf1yGPmGO5r7F8ykIdiA+ILEU/FM6iugkada0NzhO3j5o7yk+NMku
2Bd/nfRYx0Le+4iisPMvMRCZHFf6YeSZoqidiiyMyjti9xFWJMKMMFhWeSRzPfn4opp9IokK922R
S+25BKPfZhmtv095h1VFMU7xSoNqrGY6YFl25ddUPggzed27tNWDKwNse1DsNBF2yojrML5KhPKk
DqTw/Fnvz3NDDawMYrOF0w2WM4kWBczfW5aCtmNyNRkkT+2QNNdxRNlgodBD5iCbvtXEz9qCDWn/
2EmJvJvBlEuIoLu8jfq4iW1w3ovJlkFE7AsBxRubtvWAEs+q3582eRhg69PIKjcnLlFZh9VuIRYS
gk9w47BN9uYm8rBYeHKjbp1t6AUYmuPr5rhn4yiNpzaEnHRfZQFnmbAoaSRIvtNwkXsm+3zq9pbC
xaTvBg7okVZtpHrnxBpDEySDQAMv02t+KaMK+CCU2aD9LzMzseEmJrE+5Fj3a90IRoIsCPbGlIFb
+Nmc7kpgN/2BOvuLy0yxG2LcGKHejiQKCCZmjsadGHnzt9h5r1LqtZGm0hZGFyzljf6FpaRECta/
DAgG/7RtxjC0gxR0/u7at6QVIigzsImiQao8J1ibdNXqKipp+tOybeysW53SPGgIKvDs6XNQ4QsM
a+wMHKVPUa8kWNcB2d69d+StYyGQLkaRtD7PN0hdWUKptX5+a+Wy2f5F4XkF7YHzyRTtS6kGdtIJ
xZP1hHiHDpaWFvA732cH/ZR8uH4TeiP78MAs56i7/Mc8IzfNmUT5V51DWHCTTzqJ4qkxpoSboAXa
NnYEL9FkM5y+k6o4NII56xyEuXhw5WVSASugb5T8sR9d0j82uHaDMbDfJvR4cSDccsL7iG3TBNam
Gh8hpt8Qe5IZJsxh2zSfVudOEE8TiwZywnYbwrCy5Fdw34mLC0zAt6QU/T01GwgG3QtrTal7w5T8
KA37LW/3Jp50eryqH3PUCwhjSBj0iMFd2D5cHvUeG7sJvXoxAvGfKXtX+QJ6Ltka0bIkLHHflqNv
EJR9a4jjo5Wv/vn1gt0QJMPJ5McMrRF6+1vV9tX8GNkc2lplfpMhLR2BzP1FtiKzoeg+2J62NoL/
ydzGGyOecdBsXSlNEWky9gO0RHs5puTyiTrQ0PEqI5MBzXr57hLfZRlsm6YP10K/Fnfz4AchIya3
YKvUE2IPtXetrQek06eypE5nEZur97vkpJ0SC/PZSwi9FCVy5MKekM1jy3xVkeS/461/0W2gSnj1
Eb6GMHKv0qE2hyfcNVaG1RBhrfUJQATdj8I+QfIOW1WSYHN0V70+tVy99evrcH5iHOSXX6NbnELx
ngabUi2vOBST3yLSMsTS3OiRhPaZxCT5PTqIXZ1OQ6GXJckxarS26mLJopS5w9zhwBTsRAy7Tv+F
sAxkcbyDGyrggFj+FL7Bsvi7Iwxii8cTiHa6QrM7FZd1FJvVEY9KRs5rZuzkLU725bYwQN0URPQY
oFNJ3X4k51wfAIDorTp2aPg0a0XmgyrZ0PWI7+7Vt3yPBw/abIMOcTh+aFF8eJe5GZ9+v75zGXSx
aGEs5Wx9YaZIjCjiyoO2aL+tt4KdVrn0bTIhTPyu1O2w1O9qAtPYc2AZSnELyTr0qJAvQVlY3Ael
mhpBPTIyqLHICPUPnaxurlpVCxFdWmg5nOQDW4vji48SQniIZREX/XWo+4e4qlfNACz/G6sNGFZT
hdWRJe0uPJCOr+X+EK3fTXrBH1UfpYeXSvcAQLgPsCHgKLWWfn+Bs8hppRS7asDcRRDN09La8Rxe
agSL0/jSvMKizDVzTqWMeVM6tGebidC/2UvdTjStm+xQ8/W0t+rlBW7zLCce1inkCqWzOJ9oTcuG
xEcK50ckGtuYatQiE8lBqEJodn6LcOje6K6Tmrag6nKct1/u0RtUnGRq037hMh6ijIYA/NEaXZTj
BnPzNyi1o4pAQbLWBCyYbZRTJ1TTgi97i3oFMWJPH+pVd9KmLUI/cvru+E8l7FxlNgbWPOujB70L
l654lCpf7UBMtD8uYvelgmvmk40wnNSPwA7nWSPz1XLslpjaw+iGz87zBwYgE3wtGqOaYWjIJBlR
misANc57xWRJCGfGaYWo3NUvSIUUMeUcsU6vl5mngM7ZUBCY+fu+u3atMuoN5ons+Mv+jDiygWdS
Rux00v/R0Kh5Y0Vsnlb/XlSqYw4gIIkpilrpkHQHyQa9FIQ86bDl5yvIoROC4P3s+EteQlVzFkLn
iIzoYfV+DMXOs8TTcBA1yeLBV+v8lIaeX7DAOH0prA+SxXSM4hj9P6e602Chm3I6aLz49YY/5VXE
qC1LZvroF+k/0KRFzS8RLjrXMRFViIbCrC9HEneOXA47uA0lVnqf4+4mC/ss608jpZrL8/w1mI40
8CXQwopBCKkADmH+eqxNMR5im84c6KDnYNWnvg25fzXYvmeoB6d1zqmnb/V+4dZBhzJXYqJwuyAJ
wzCCdb34Xq1RGMWWDPoKYkIuUQOvcQ3rHYmRxaHFfnllAVByt/slYFvQeB+j7I77EC2/kzUmgmEL
t5KAPE7UefFs6Csl0cwzNNPU1s55bq8gpBASg0xeawCdvaM56b3+wQH7M/z+v0Yl7JPgu8ehKdcR
vTJpeWlgKMoJjTd4A4y0wGjoQQ0S8rzAs2b90dceJY5YUUu9atUzo8NsYYMZ571sLiSOsswGSQXs
Z0TlPOemxudgEoyuYH4B6i39KpXEwXKORPBC/5o+vrMRgGZhqXFF9Acym2MSTPvSDOJ2Pssnl8KL
IlG8wARVat/alcHehN5bXtYlCDpkPcxuCIQzfLrG3U95Kd6KtXmNWrKBBFu49d8zIjUu/8NCfFKY
7rVNGTcYtpSGPGIF1sxRJEuHm66EWcL8S1UA8ceBeQe0BFFnuvTfXjTT6NUTNnJ9nRAzSaJdI6PU
BcLkKhznKfdZxJe6wY0l8LG+ECIETBzznCc2wUtoP+wY/n3B3lcxWfZ9G6VhD3iXqKaQltkii7MD
wHVgA1v6+LRrBWSTIudgfkPDDvTUWANa/5I6sPt3BNJ5ltHHJPm+b5ttE2NQIrT5OZMT56LYQOmO
utpYFu1HH3K6oDaStjHojYIizlYAHT0zP01SkfeUAvjetyUkYViiQUKMOGaGBDZOAnxE+XMR5VWl
3SZJqUtrKTSAloxCZYU0eEq8CVSLjSCdG1eqjVzv2grf14MwbT6x2hUiKjyumNNfCK9RBaivylJm
v/mOhu7ns8Z+zIT5FwQN6G383Lt4S3UFSG8cEBpttVxi9Vc60n72a7iuQUNg7xX3/vzH0mzodH/z
yueSCRigzeMqj1YfNoRleEB21Z+Sk9HHlPCsoYy3ZFm4CI9U97xpxkYw3HHVxXGEciKgVXn3fdP+
9JQL1EoJOWCWtDSUhdp/IX3UbSTUopkrF6v/EkUsLepTGes9aYHXf8EsCGHqmHYyv8ehBcbtigoW
f1XLGuYm47hOSEXLdOqSAxLpSxwIwNxuM3mXQsTEzIg0UAEYrrsrpO7bfSW6MgnsZF3fyaApb1q1
Nu4JybE2miaDV6YSAVPHC2YGh6IUwwE+4InobLmvjo+wYFlsmwbU8lPmThhYzbDwbvMdOd1uU+mW
j1BnGGAAWd6J5halkP/UPwiDslz6QVt7f6mG4i+x2NG4cU1AFeTTKJEkKhUHyUIiDNXLSa6ITqd2
9Hdgqonfpnz7zFSaPp3C0oJxsTdvSpjr2swc5kAF7tU2n6dWPAAnlaxw/I6oPfGgdvMEgfKCec8C
hl2FZBFQhWeJGykQU3H/Pb7m/l2BuTPwd96Znif3QudE8yFbPVi0lPy9nxoSUeNSn32g6wu5VI32
izuCoTG5qhtyKAdVuQf9etcLZoIw7T3zVZuzmUl0rRI+TOdG4eYvZW+tH9sJswwlfwuc5dwjsvnU
5GFNH/Su5d2NyymXjk6V2LCw3M4edRrsjZkAhG1lN4zUWBw5MXXQdlN4b6JWF1NNBkAeAR+Az5TA
EXK1IqTdi3UfgHjTvUDiUWWOJXdv5DOezw6yc3++dPGUkmVOBY1TZ7Yz418tGspbsaW1dL3Y8X5b
EDvllxbSQuWMADUtIwcbsi/qRlHvqygmMX2Hdkn/ZbtwLCYki6cJm1kgTrfpqO43HoK6xtzsoTz/
xjDqfiE+FIRtBzdQOW/qrxEvzKAOyKBxNKp/NI1UmTxTRgrF/31HROjUPsDOwubp9ZEFPWOiuaqQ
MY0xNE66bMRnY3Vk2hzSXGy+q5QtMcdQxTZPTd+O5gJb/kHx0mYU+GdD99E1N6fGM2PfuFD41/LT
cTfs39RJiimK2q2WOtX3xG/EJRqmEWGu8Z5qzkqXvExYIo25jm5FBt9yt1QDwiTjgPcr2S/QQ6m5
87icFxLFefzH7EsHD0WYLMKPdrz2O0K7RTEG4iuJuDhzLP5J1+ucUIFKojAhKPq8J1cNvTm/jvB3
ZAoUWOU6glnzWJM3pXQ3BfJizuGMcjNjqhFN1wCoTeN56XH7a4Jeo/2elznpUex03dXE1DpNIEbv
4E+k1qQ3Pd9z5kxvfZyvEZimio9b6RdXBDpvA6axi+H7fZ31J0QcIlyLEgGWiRt8vUJobLuJ/sME
KDB277twSIDNA22TjKyOhLRCm6x+hZUwWw6rl+3jIASn7SlIKMnEnJiM2MgmtqGnstfPSuNv9GVV
4IcsAhGTHnk3Wk/xBWYQ47CzVu0R0KUeIw1B5ogjcXhlCv1LLiYfmVryIWZpbFobvZ9rTO3U7M24
QwMe6cjYgaFgFx9DJhlQxDlbp4iq1kYDSl2k57Uwo6PFoeRDBYKYNokazbhjNQ4K/0UvqMaY1iCP
ng2jvTXyQf2+sJ5g8KdddquCcg+HuEzDOcrU1UvsnnVRMX3CZhMqT5WcBnybyH9wcUI9XlBXHflx
2QhIswdWvc4LqFSVS+VRd2kQcp/laPBvfloVJa4pO4qd9U/ogC7DjeGnCW9v7oi7uFbHJe5YCdGu
5ZD1+ojsTUfx11+H9F1gwzXyGG8Ps/r/F8A7MXBkaQ60quXTZJHLh80/avtLW4uspxg9K3HUOHBy
K8eLqyd1xmZTGfjP7zK+LnX1VTEolD8gUNptWU0suJ4viab/3X30aKE5GKWZTJAoJKEKpjWPvdq4
+xnSJ+TbOjmTJtwBCYIbdWNGlBcw4PkT/qVlUgaXLpqrGnjOd3kBk6agF4kPp6BfboeTzUCnFQCK
GIUqkZZgdv1DvrLt+jRn6XZMsEzeIScg5rRjgu01uXga9NV+OmYG1H0KD5VUCmjCi95SToCtnxyf
pNuJUMTRSG4NgktXK6KxpDkCsE7kGuleg61+wg15CLjZizborPJVn//zwL96ir1AHkk5BtFrokXi
h3RChmRUYQPe9lW0+eBYHC/qJzUehYgfE66kSHcLRk5TUVqyQg8GPYLcN6PM8Y6faoFrSp0WQvto
qRGJzBQJLnGu6LeUGdYUPqoCMhGTmX0mlOoPFX8NrvwFHWgY0f5kTHdcsJc3HJwEF3ij+1oRLS0b
W5rVBbmJmj0SVWEBVDzAdpQOcp5bFqAbbCEpBFCYtyz1ruiCiL4YPqrKCjrR24+hXoGd6Ag7+iS9
rG737Itw/hedwipU8hN/U/llq47Xt4iJwX3BXeRwKt9csQY1E6oPN7YDOu2a2QjAojhcXkCUKe62
1zYhReojOZ29VnTAhvAEcm5ZcHtn0F0T3QD0U1VqbLwTjD8oDm3iTS9Nto3mApd9kDwPxh9a52tn
psL5jbhCLB05CMqi5L+FjFXCmOTaij4uiES4IXGQMRn/Fg9yFOw4ADF47fZPgXLsbFxYvFNVDZ+O
dqslaqPwn4mU5XezlJKrNMBo1Uk0rG8GlP7T4JcbxjeAtQ6zt+dgh6Z9aDeLcxBfMQ4IBEpt+WQP
Zn7x0ymbSirv6Z2NUyB+/xTbbHwhzY7GC1t/348qUA3RfhOKxgweC1AmrmXhvqo8AkgZLgpFynlh
r/nUt1jkQczt51gnkMHDguWnXXqD1lcLmEP0ZsLb9CFs/nwMOqA47lSnp80ruHWAKixb3EQn/NUz
iK0gDIA87Mipc3jddZm+n7lScR4iPhx5ETGPZay/nSkAxjlW56KGhOdJkAdUfCEAj6W3rGYbmHir
2y5WLY1Sw/LSmFltZwqgxR7DXeE9NU2dCq2tnE+b5SlmaVHmCM+St3aEZgcyZDGkMOJPlWRHoniN
FBHYoZnbvVouLpP8CwR4Z09qHILd5k7pC2kEKdFa27SHz+l+Hf77sqiYeY+YMm/z5JS8J1mxunOx
TWXClghXD/+DaaELOSyCg0WZKOmcqyt3PPHNh+0DgMvVSOY93KB36Ownnzz3m9GYXVbIAEo6iDSl
i8ReirvsTKiufb8HvIf1UI4MhU44Qbq/zxyDmcQF5gdr7aq18BbWYpQQrzPGY+axMJEjCEL/a5Db
Ed8hNljtjJLIFSbL5LyGcAMmaX9oANmDiCOPNT8bny/2y+rNwhdc/BE3BLhjWuShnhZBQzJVCWmZ
PvVozuBLx48GWCC+z2SA2yv7lRMVVW4IMaiJYpigp65AIWfyGVy3eu4uMha/yszkWxborpmT9Mdj
wYqGeqXChCxZTkEymgQ+M/PhPPLUisXTBNbk1J35qOF0zNl2ZFD+MZk7gqlfOlzCPlVUr3iXMF/V
6/QdPNgoMR4RLAu7svV+T+L/XuAiHsrQk12gToJmkzIQLq6yVOW2HLJDD4G3eW1CHNIz8DIqOm2K
lJiEYkYlOCOJquFAGF1q7ZWvBVfekZBAcfYFz2uw2fETrktTcywPt6TucozEz7ycf5Fn0KZ1O6i3
Qbx5ZdWzy5rJcWIl6O29WCoyCIAVprkcFt5ZJ2uDhjzGlcNBVKks/t60448N55bkT4wVsGHkY5po
AlTSxDNnSG2bfu0prHZtqUAjzCwCyMUGu5Ny2gPnjtnzkWljswW772Op7ODEGPD1+uMWV+uJh3Tl
Ah/poflJ4sa5sTj+0AZh7XO7CNEc+jS6u7MRiVijb3lFvuts0yYIke2Ho6f7ke7jSLP/Ege3oNnN
VYjsQv7//0995wDZw6VpRT/mYtsyPzZo4Ci8pb/Gs28zEcPMsbyzNkd0K7s5NXs3JntDaZVH+MVK
X/vu7muO1Jns/JWAsTe1J9ny5C4dOEUHewy4qWqODNUvBbLuD8jUFyWn6t2dtkVkiLnrsYs+0cQD
K60Ukug1f+9rZh1gfKlWwZfiZNnPiPn4BglHhSLcgxF80b76Imlzth+oztaTmbCInR/tDDJdjFHl
/GdvoiJp61Mk54QGzk0x6jjQRDrwPRaTyLQkGPMra2oGMRgitEb+jy5XJcQGCRFbQ1qh5Se8KNg5
lM7o5Z9ga7mdyaZ/QxHvO3tpr3KZVEQ/j79VUE4AvIfd5/F0OLvO11Ve5zdjpR+yMnPwqJzLoZpm
UMmdIxS8UNtHHfgfqACkipty7/0gzyMP3mEcfbpWbyzErvT6wsXiuodcHwU6dCnugRdRjJ/KLqUD
WOMAT9cU6MAbK66VbIPyDfL4HQKgF9etXHuocBWf0KsHDAvqvh/9yqbiOcA8eY0kJUPSQdwCQqpI
WToCuA7K69xv8fwZ+CCK0Lc90Vyoslf1H2BxocuzWIcWKLlPgY3XFFsLqZK72ycZv8UIj6KxBloj
y+K2G1rRTwiz43r5eIU++JNVV3ztFaAYfX1LZfaYbGJ5/WQ1GmP1wemYErq+Ps0k4/ojcJ9402EN
IbK41TujIkZ5vLnQ0BbaAcGNOB9KGrOiBbPPXarzoZ4Xa37qoffGlP68mE59doaJa9rU0WQ8sQnX
jPH4CvPsSGr/nBqQ7+jQtezxVtq2lIOZTeVSSh+UseQl5fdUfhgoCa7LN8ykc4XCpQ7bd30BLh5g
TzA0Xh6rIDqRMoSr17D0/kr99hNvRoJNAExtHTYT57MOF0poUbN0dHrsDQ6thIJMnFDT73faAHF4
zb/MSyXo54uAJL2sY72QXYNb64Tsb8ex4q/6uz/IMhZekYuvcBK1padQg5buvQjIwIzevgG+MzDz
qyaJoWuvsGIpAlmc4I7076TDPZ58HG6VzB7prWr1k5t82qRbt/370iEo7N+mn/qMZYLarmn8XICT
3mEXhwA2vK770KjFuaHiQbcVCHPIYNME+433pQb8rQJqdwCtkM8Sw3eprVREDFmrAf2zT8PwJcvL
zk1KSvfyoJXGWcNmnDij3vWmsnp7R1Ei4TvX9/vQykruO0ZBLt/EmfgKlPoIxJ2b3byYTJjFVdbo
DuvuYHNdQvys84tfWUkiPD1L2eueJ2FgTwu2REQCdATHJoIh17+xY87d3A5W575xft3pMnbeN4B2
JXO8OCbNf2oJn9lWprrcw0TVWQf0VKWODFdGHEZA0EmLpqYmpQW88r1FhhvHB0tU8+0TCMIPR9kY
16DvP27TVdIFbt9Pe/o5CUDc2EuaRBJniMXltCflbBAp71KjfP4lhp9hav7GEnp3LUqW1DUX7oJU
3U+KSIJQoxjtthPFTHheh9N/leRG+8HwR7mY/VZPcabIAoSfpkTpZHUtPoy0KpdpL+/lg0mhflFT
al2iQ+maBbxei8RLsrB3hk6/I24HYiDYslXpova0WtG/LEM75h+NUvCqhTz9BtxxVXyXHZYU1/kD
YsANPQ/J68+5dSRQldKZgtR9/UmnGtmiYNzaqU00vIwpNhC1Big3Emfr/GdoRZZ17AU17SFMEv9W
6csk/x3KETNFAhatY8G7LqsTaJBz0cG7xx4G5VyfEHrUXijKHZi9PBgS/hVjwyi7ZvBxz4+7q7lq
SD6RREhonpH7WIwNN5kr3rupWwt2CuOM6LmpUj82jd+QAgRGw9+seIKJ6f5lSb31YoSZWAMBWrvb
YF8V9JxjjVa8hMu0WF+oLncISTWE2vaIJVJlf7wkat1Wxv/WzVJBMx7GLMyeYgtfoeE2CSqEPrFA
RgDxFN/kzFEYcOWVpCYUTnG7cRs81CMQwFjnvqwCAIcPzH+F1ZC9kmpZ1LEubM4zAM4bFD41V54n
oQA/6qaMkzo/oNHZlBtIElkXokO2VkZO3zziVHETOWA02VPVxy4iad8JaB6PoO/RyWRYB8uzrZ8D
YczgezVXO1lHCIJVCWz/vskZZRZygRFTolPD6ZZGLYKDPxzC0Qlerb7V+6G91btswHBqLAcZWvzt
i6sZrSd/7TqbvKvSwgTaJHagiQRTw/xs5akKzDFFOrOvdfecW/RSUrVPUQcGcOHwgmlfzA1PzBhC
1IjrSUN02EwEk1ZUSafUPfSeqpLRBwDK9uXWL8OxIp1FGxKGbD2tlSP5JPrGjI2LoiVzOxf18OnO
fsA3pi6x/hpB2jd17i59ClPoi/bG7O1t9V33UXOpbsN/ca2NtRsA1RBj+1PhtM346j1gnuKDDxqY
vI7maBqF6gIbGuue7s62nGBKTf39Aj1bpZ7dgfUcN23SL684jdHHbou6FBOIXzNDB1Ymg6bOSndE
2XYYhOrWXol7kbWnzoEIzYGpP6o5MYNgyrFmklGkGaqRLERQwax/EFSvtypqFjUoQ5Q8Tr9KcHVR
qO6T6qW2iOmllIlmDxr1lOQmWEp8tT+MK5/L6STCWM7llIQkk1BmFDrcDmAyB+57b3KNm7JPw4jt
HfuYPCtwkO6sEwQNoAmq0e8FhQV4gwfyz2JtqOAewI1hvKtAMwFc/P4pOI++LAZbY90Vt1p3q/AF
RoQuWjtVN833l78u6qGl/IRWGGAJepBuj6HodA99t2SGDxuCUDq43t9s5sfeIv1NTBopV2VtO+pL
RxaTYrEeXwcH7tmu39k0K+0OSHf2qEftTmvlOgAefKwPFbuYb/T/tQXn0Boi6dw+hBX3z5zd3xvp
YiwLsVpFRcJ4wKpSOhgqc1JLy3nCjAK3DomBmwdKvG5PshDH9EATRLxVfq2yFAh0IBUjqvaEuoxD
6jQMtY8RpJzSzoL4QMbTs3b2QoIfLy9AbqMvlxFqlkRoqUE63ZTYDOf1hExk4T+xIH+E3eGoLVSs
Y0vMEdfQBENsfai7sOauGSOpRafcMHautA3HaWUc/1jtL+hPWQW29FNb37ngBZbU6qZM9H8x2aal
VV6Ph8zCn/l7Gh644UMrF37D664LW/uCkc6b+aWC2n3Y12OMjz7HV1RntudHlb0bvE5Ee0oeodkK
xKtYGTo71ZnUHSo7hOothXsganQRtC9YzDyoqHUK7PYYe40SbcCyC/uVTLXlKgYGLY+Cl92t+LS8
u2lhFOcwS+InCll/QMyxGU4hsTc4Fn9y19L8qtS8ovHwjALew33463cyAH9bnq6uZzEQ5nr9+UAr
q5gOphefVnEnKEftcdONIDoPGdMWJwLhTEOy2668WO4aUru8BD3x9KF8sH9zPDDV96SFJG8gV320
tRiomO4EoYMXSe7EzomSMkpQiIAOnNarAW0wbTitSL0g5uFcji3KdjgqOvZRr8aJIkJtGXMTFbkf
fgrqpGefOOrdmnnrBzFtTi1oXS+TEOQw7LE261dRAZnJl+cAwSF0C6sbeiG26v5cV9ibisoJjxHX
/USUl6RqlJWIDoYzWAMJrAwfpPP01o3cz0J/zc4T+Pc0EkfWXlxjcaXOuxew/JqncTpBLBdp9F/U
aR52yUb4y7cYDbDzP4BG5GAU2dn6g9C7XLYJkkVDQIHNfst/L1+etTnuKr1dJ24fJQQ35IhLxdtj
IGi46C3ovy56tMDMFuCF6yomujO6ObsLHQR2QmKvdb6d/xYWgW8w/4ied1YBobMH2qts+0LFqtau
JH6BQWHPVp8ymgwL8D+h1MzUUtObqSL+Bk2PZzI/WIUl03a6dZmcvxw942QekPF/Ixm55hPsnyCg
f9M5XCGhy2fYsXMDGMQL+u0o/hQACQC3zyuhHjf5V7hiJXdptVKjzxkBU/2+0EM95rtvT/yJvphw
wn4bKSGXRGJBdNqCtqHMQ+KFm6zq6vWNWQudGolETNW3WmZEusU0ZOJT5E4ddhempXSuJLVOP/dZ
ZeRIIfIeh/r8B7sTxzLvFFbTwTPDLcS4Dqhm20n8cZkXSwRYrmXHyqAuMz64vMDYbWVB5Omz9vgz
vBGGW369hkkUSgxr1Kiftob1/N9f7k2fQlo9/wJjdzOU6hJTi8mvFZtBTk5zFEMf80hzoSnO2fmJ
ChWvB4A/8YOYmFaTucTS0HVaupjXKlPOP40Jq1pfydfc+nASg/p7nHoPj9vMEc7Lo1hI/lhv1UJc
Qh14XYvuPgSyDW/Fbh+tPhRjzf5fR/8XadTMI9Vxk2wkoBGKrDua0VQBx32xaEvF59wFfciH6bNf
aHg3PxbFfagD8a5x/VuKkQksTHk5SikQmFgd0kEAEof08MoDnQu79X+vOJftV1GLzObtk0cHKG0w
xK+uIw76oAOzforU179YNkWdG+wWxmwktNRGd4FIyNpIDrSC8bF/XRwDUiu+18Er7u7NywTCDAoO
c16Tt77W/5N0QjQQcEMI4mKnIj7luxjmLOFwv5o4bn9kfKzOb8NDa+UB6DvrHMvE/0ksXVA11B1g
a3wuuaWwFqBuzgtQDC5S49HtlxPYYWPwgBP3b3/Qolmke/mB6GTQdnL3YD+M5d43QBB9VkPvBpWE
bYbvHVZ4T/Fot47ghxqiJKrRQq7YgvVs+d4jewTYPzNwBz/hIO/dSA+a3JEllcn35GPvr9UWiIvo
BbxJHnUFrVPicaO6O4Sbul/dMLT0FsShiCwhgtoM3+N6dM7Ez4gFS1hjbHRLtxfgBp/U/prbp+Ht
Naa8JSIDsQWGPA5anv41fY3lrMTjSdJTfuj7TWAaHJE4OEpMile0y8rWs1plf4SFCaBQpV5dxOBh
7B6CL5siUJLsfwCCOhUXPelzU60sibWSHF1Vi5KwHuUULLsBZ5rVuveAo3NsioqGK+E2OjRE/RJp
TtP9dE8CSVBe7IcuiQD5LroGp0bOa8n2K4ZJJNX3PJ6tRkXyUEa4CVnPKulyQbZb0R2Y54yhfmDK
JCX1l3a/9EB/KydEYFE53znR81eisuxxvh8wyKZiFknJX2cX0q15vuWsiv2kz+mtg9Ce60WHCpP2
C9GItBX/H8n15IHL3m7GA0Gtsj6DoXNpKihTFUFP2HA6sh1qNizXE6VQ+kZ592idDf4cO3vYjnDE
2cPDUg515PcHXLAmJI+p1HroV7a+sxJ+84cAhIEQ7REBICRpupuwyKIoD7vTu253rKSUAo9RHQAg
2yQjXYqofvM9YJkRe9f6WnWX+SgOFXK96l+7qUPKpupubNpCRWCgEdm2w1GjnWOdvTmtdadw2FQv
nkCMEvSASjNa0uhXOzoc+l0lXE4sTijABu77d2WTUmpoEkyzsehbKbVi+ZOdbKNMkvK7G8gntkKS
ZT0K3hZ7gY6bVIgLEwYApJ3J6fWAwPL7sl3cm2rBGQUKq18XxHtkTmRuU3UhsyTJT4De004C/zV1
gopJGaKncVmLZGyBSXdlNGHosZ6ff98RFHKfTBew93KUZj8a62eEnqzCljWxaEiAFV527tQWlO6V
4AcpiC8COG4AoXYBEHsWQrizSN/INJnLlT6TAlLlllQn6sLSU8xzTD4hE50Nr3EBrdfPU/j9n5Wm
bNy7/LR6GASN1Q0qDyxtWbSF3nRLg6bRiGhhmc5h+GxXCFftuOrgYu8gBeThN/D7ExnLmFrVpJ/8
Iyv981BEu8ZR0FdPJ+OAU35yy5p3fSpCBeIOgeRMYD/S6gIGKPgBtDMAQRVyURbJGesffAJuLDae
ky2J4Lzv01dG0uL+xiPlqls9QbM5o3LFqpwScdB1Hhuxpxd36jrng//U8BOnc1xz/E4t4S7oFoEv
4naqhb/mi4TEhIVrFw6Wlam2MPEjnQA5XJ59PN63zppBwiyvXCugFHvxTIKCJk82rpV6m46P38NR
EZzxnEDxqCnPFN85AgVawMVrelKGTNQ0v4SJutek7/ti3gxbupEPOdzR8Jl8lVQLyJs7ySNeRAX8
2d5wKaQdW+PeWqDOUVpEoetdUQVn93NzXzG/MMKphJJa3mO8Fy4Arp/fhJ5rNVEYFyDA/syTwFzh
gO/QEofySuBEKWi+AkyOaudKgUgYAm0zApM/fwCMXSwuHnkDsVuYeYbBCa5FRrocYPJK6HqDc+pu
93XeJFiMljzwTK/9ejITx52gkBdWT0WnX8lS7WW7GL+vNtnG/b1EFMHTD3rM/BZN49XUzdKTkI9i
0+7jDdcRIaFFzbwDjaEkSTlS1UE9/CfMvQnzV021yzecu1X2w5qyXfEI4p7B+ouDrbgxHF6kRigv
tm0UNFMIdlgqjP9Byr5cUpHjcVRRNqbV7Gpyytbb2fASJlecPQdOsXqftquUvkHbHLfpDeOT7XRQ
QXPmfP74myyi1l/qF7K2PFYzWKqWDOCwJfiPMqG4VNMEb1AxoNIMh7ioQvoIUDilA6FKXpFx3BSk
TvzRhNPGYoN5c2GF9zhqQ2nmw+EbQmeoXAOd7cYE5ozhax1o0mw9Cp2q2nNSSiWm2GLRI7/0ojFC
nXTb9nau37yDGcK3rXgUZ7xtwnF5M0CEdgP7GbAesPg1z25M3gsfNe51ot46gJp9HyJpawYxvYGX
fZADMiJmhhOJaqsjo6AXThQwT+cpuDk2VtNPMeMnInmd95qvmZuUND6p54/ydJc4RqXBrteVTqE9
R6B0ReTd3EdW91gYjLu5I3K+7XqYn7lR8fh8BmRmR8FDrOpcYhXhGG6u8aOm9XxC1QoteOFjrsFX
tMyHZGomOjHjdyS0uFn/3U93xdD0/qPnJf9fdXVPagRL2iL1+lwgm4LxOdGbstHrZ4qN6VewabRj
2ALmBjQ+8oc6c3kq5ypr3ZrE19lFh1jG2rfZRP8aEBKn8Q/ZFOF3ULtlOo+sfRgzOcjTNScaEXig
SC7yWQ3UM2MtaDDeF2lzYfXi4s28YKbe7EBIPRBTq5GnqfPbJBx414Z+sRWP2JsFePboRJH57d9H
gEGnu31Hi0bdqn1tzD8JjFQP/DB9N189zFkaBNlHrtebgab61eo5J17cwm3j12IvUIph3gdXY5La
SfE0rl/j9TLnqXvAg0/xlLpkX9Y6l9nnj2au4eCriVwV1n4F2CSbaPMG9Cu8h85QDp5g0JKzzsi+
juijTsTxsI4Vio6qf9MW4U8ypYw81AeCkxw7TFy3QdldS4zkCmBDfe7OutFvGFtPXQxAYGz/doCs
1j5InfoP16BwhGMozarhpAqiakAT4ElGmvd08ujb/YLGGPjpp35kPRcyu5keBH8V6okSEPyxT7Ok
dCbEi69XnqPwRS9/WEuro6sChsRS86NkTLqaNLJOah4JYVXWl0E2GvB4f4kBojeQjYoMGXrpIqLX
HG4eAQScY14/1NuCLVGfoOcOEjuwEwDrZf6vCfLTOy6XOA+o78LtA2XTpMC07NgpUgqOv3nZ1PA9
chTzpbglRgnAMrFuAs322PvZk8oWTECl3Y+vw1htLOSGqIWkS85r5aGAJXVHjmnuPk5iUaD43OhU
iuvObo6GH1ekLUbEl8V6EYKXT/NlVJxWFTR0UOP8ZkStAdZZ5r2XgLN1BdiJUXrPYf3pnax8OtoD
zr1NzwG5i4LPseO4seczymMsVO1kfM/ivPPK9U0NGHf9Y4qOD7+LGvL1P4oCRSO4+wsD83VtWex2
Hd5OHe5cp9Uhsub9YLavgWNoiz4QUHuTniheS4cDRHoPEt04lsIqoSTuGmzg8kkNi+qoPfKkt13W
L5YmikowWRWWYeuRc7/DcKg28DnQcMhA3sq2omO092lHeCeeajwW+ryht3e2TBZMKbvP39m6NwQa
2QK6rNKoCla92SYCJbzpThQKOt19ftklWJIVcw+7D6RGJfovPfMxW7+V0Qxe4QeC27CRVk/SC+PR
ohtAFkUT+/vUc29vS4bEXmXAYXowSiU4IH/1HcKCFF+fFixY7jpejbF13YekQ2M7DaFOyHPc2BU1
x6PFfDSJ6iArHuf4M1+N6N88aCGEFMqtnuFdmgnEFwA+H5ZIW5bnJOAsmHTf0gJ35NKYeScHChP7
tILQBqUK9ckQMO+Lz1loIlg7vpjW9o/gf73tP1Y+KZQNVoMVcNMxpOiiAUdqTFwxPYAhYliezGbj
e0q5OG0fzoA7NdZCR60ssjbgu0xyvMpVAcZ5aA0Xng+gsVqWcZTY+YWzYf+DAtN8NeUgpENhs9xO
J7Y3djFKjzAWy62wIPHcmd6CjuOM0qG7xrFCNoogUUFSzBy0PzuHC5Q3L2JzK8ooSbBXOOo1AyoB
f/V2+r3ODcj4gxg0Sjw/ekKBU30qtNapF15xTKV6DOVKeOBHl3RgufI0RenkwiJ65Dluy3h1wS6h
25Sg4QfyD4Nypyo/zOA6ga9ef58CZhNn4VnCCGtjmMMLocLLquQ+TTgtux9pJ+s+25M+eZSuL2Yq
FX6ROtrEztAejVuuFgzDnfWiSL2KkVXYC7WxQ/5nv/v/GNo5hb136WQRwqcTmk2hqnNJ0vPamdym
OM0u5sKOgrinGIm+i4DJ3yCz9lmQDOGBL3iTbgWC5XDEat3Qs4t+TrhrRNlXYHt/dGa4jD22RFlk
Vs0RY9uHFK1KjRaIlV8EOTZl1PjkPEpNDg5/Mcox1wb5FtmQdDI0kge+eBkw2ykH3SXe4l8YOpQz
RIgdw8TmDzrb5+sG5s56+VqaFQfYFQb2wN7ORUxQqFacS0SZfGZN39ZalYoQWO4zkCKE3VbdVXK2
7aeR8BZiK1f295RuX41wx+fPg/+I/BjrKoHu8lQ1fcwjStGmbQtWS4uGlIjX1RZBv0F7lk0765xp
tYM+bpgL6gHES+BWTwvaMY6lcdMZJ7ATpK/UaZEe/EX29hM3XsuTlZApqp9EnIQztcHy+PqXAvyf
ZMUMHqCpQAoGYgJs1tP0Nzsb85ADELAtP+ThEp5taLb3BEdvLVDYJ8Tj/Tn5lUk606iJnbM9y9v3
LLwm2ftmEPibmOlpqxFzxv+W1Vx9j+gHmmVcsUlwjbfZ9/1LinyOPcVn7W9E/cZ49ZgKuGcKt3xq
ZoeoMre6ORMQG2n3qted7l6q7omMD5GDajMMXoom3ejIoLm4Ps5+mrvkzRaCYNV4ap3KnyI7ssuB
Vmgbk3q9N/SB3RJXXexm5BRNGBwWlRdsLwqvCOjZ3787UTT2mScipL6tTd7zQ8dzzSdFdrR5V/oz
lkVmh/+oK17CKMCTFT+CX1Wt2Ray76S6p2p2nnEL9ZwD+rM+8kDMw6tXPY1QEP9brIwWQHlIVSqL
wRxPozMLoA0Afr5El2NaFJr8nbSsnSMG0gCs00/raUYZFhLZ2cNe+/mQEdLUctqbSxxKNmK3hBzc
VsXoEmLGvk/oXWebM1/JEot+sq6wniBpm6HcdGG0i4V1mE+yqVUJvo9+Sc9H2RQiVNxQFXEn09F+
PADxbiQjkJWlQ+U1X4j6EXxlwgUj0L5wGX2FSK/0BIC9GyoVuvSqONWdtsIbsR8OzPLbQv/7c+vx
GAqMLyHaDBTJrhZyAUrwno8TcXx8eowNF34aU/NPsem2vVhvXtOBnj83snBKapnz+lVlPKteK0ki
QW2n7Scng73yLCK7Xiv4O+RKOkC+/TJiWL50ADOb56Do5Vp3ZBOfaVJ01Vk7y8KmsSFd2lmQrE2q
3ziwyPYZzy5tUg0mMV9V9H6bZYDlkGPxtL1WQ72InFOQo8YiLgP95Gjp0YoRy68WShtSAgSiW3Vu
cOHz4kIFjyKJgkWNTcrFDE70kFJFH2mgBfYyxxGzZYm/Zq2ws3qDFAHN1r09ouK9f2svelI+zDj5
DRKEifJESHT4sN5K/EW5vce3nXCsH0ImpffZBbxoc0g+hHTGsHvykjAzDWhMZM1Ylcyjf4bQ4483
rZ1mNwmwwZnZEY7oUzWGCAtnvISpM+my0zcpSQOQlSlGKfOY4zEiDEGo2yB35tpyQnSJYi9H6pCk
wEciFcNeWCniRBJNZmQAy1Z2K4RkkzmJj5MZtI+Q6xLvm6jak+Qj40BuQtTZ46IUf0qrcx457U9F
mea3l1zF6PKfbObO5AqjpP0Wm0SoStFb6uJjOWXfmJPWGUZErOpprwsclXfH1VIGmKVhlIJgxjHk
/4dwPcChAjLm2VPGec2ZhtzAtLQ7tOp6Kt3vS+1J22istzG0YN/Db3GKfl8z7rYIQrH68ulBSYMm
/H48uZWh8LrBXf87aJ/IKeUK9OVOx0d6YhjrEn+CvtazF5EBZuPs5Kj3XFZKc+9S9L4c999JoRIy
Re3rHuCSZaVV+1NRb4Cj9Y0bKAiwnArrALfbuQdhgCLNONNVPTa6ZxO8YvyXGIC0woPqLpCtgVHe
Y5dONI9H10m6JwS3biwlXoGZP76Cter8J6pwHdQS5vWO1NJvACx9xC7V7ckF7G2zHTAAvMWlJrwj
HIX127r/puEcr9smsk447u9zYuDxM8ltg2Hpq1KAViSMFaTBeVXW6VPduKZ1e8jSTB8KNoWzJO6b
o/t32gFkxPLmaUrHcqkm7J+uqemoabqoJY7pCt/+SxaHHlF2D75IobVLzECEHcW2VSeauVm52tAZ
JBqnEWUCrWh1WvzAI8umkYZwBgqcZRAU0dfIoHexKIofMAZuKS07TcCyuvngP6pUlm3WKaOtLJ2W
zJk0yWgDI3abrqJquQYcSR8e4Wym2s5r0ARnMXea3EO+9LohV2vnYO6Chnt+/zsKBL7Ba28V9ZB1
PEgcmh8JWyx79ZqnFnSLIqOEgSFaPZ5kzhbJ/wdo5vDqVGkp63oweDSX2sCiTS/zXv7xvrKyNM7F
dAmfAW4bL9beu5tsBB0fc1Ufl5BPDZUvc5vq8BXIVXs4z+VWdnZXRZa56wnOxuUeEBrxcTlJ4Df1
iN4jPbQWsPpsoK0kOPP7XpOoDB2YKxqR5IuL9/et485bGQ/laJOC+SY/Hx+bnTNLNEMmXLpXl1mn
UFghYSBHmaqH9icU4Z854yAFMNxImgAIPzLLyeThyemQoGQhPAmn/Pxds7isU4kpEr8lJCZ+tZGd
Ek+TX9WLTTChoX4YgyxtuQ1Rv42Tq1WyBNCaD0uYf8mc9xstUbH++fZPtQHkbQcH+a+NrwbqLHJM
1+1ahnCE9gO8exlcxQZRFqfHa/RwbiQSFRYGWC3HtlBJcvlnchoS8kHN5lMlFDb27Nfw/uUr+ur4
Cr1fMMg4Wir8oTmYjeR1yXd/LJDe/dN2qNxDdkAfYpTpqK2U9UB7dxfW42uMwao9dMFyUzFB1EsA
AzcTXeZCdB2XTfxt49FuUAUuJ8NlKfjlG3vYWxVMlnXyhRZORXfuMXWK6lPB9WOQ9LP/yT/240Qh
os+H87hM9vLAZ7Ao4kzicPl0lrFLzhlBwroeJSTNMbcMAxsxt9IowEGTqe+YZHk0AmiqAJLFxo7l
UOt+7lfmmxaVGStI1kL0KarQL1q1W219sxcQQPKtlh7A5Rld3xKDVEhHjzDU2yT/2MRycEXWrIWR
w4uce08hBPQ+M7EB76aqvL2ibyIHyzRdiKUyfoqvU+M0fiEjfeH3uCxT1s/ljQictmMF/M3zeqQY
yEPDRXQaS6Ufqp0xjzYxijx11092frTas1Em7UqV38ta6CH4NVOzWb6T+77I9mda+6dhCLs6WGCQ
CXkxF1jB6wpT2vRiJWbqbxbxZGB0V1ME/LwXOwn/5XJpYH5v6Ks7Tkqde4Qt02+cGAkZg3PfKkUi
5gfTTkIFzt9G+z+0+rhlyKDLSKmTZupRBGsFYetDMcNI+oXewjglqf8t1Zgn3RXaInLN0oE0AQqF
kvnhg0Q57c8SJ9IKL0f82jJf70FafX0r2MMf+raXBvNuYIO5pCWTtAcDNL9nVyQdwXWqXJIVkAF+
dJ7/BC4T0Q+rsjlUwfXXq/LIjpdJ9Z2T/vN22WNJ7O1WhxFmt2pqs8tdue7Y1vQaTDoXJ9d8V4t1
IXESHenLAOQwEDhEnUpjvSn+zojv01KCh/cEkGugFfDnsZ9obK+fw/RrsB60a7kKluxGJDR9HH9A
4/v68IKbupE44LOyvXDIlZVw4STUWdA/f/wv/PDoT9yV8v28k6D9bSkjmfbsuUzKE6Dn7lYDeakK
qjzJRaAvVDgq0m/x1kk9E8CKfY8vvDo8WpQej6jhCXI6RE4Kk+sRmeGSFcbS7n3MKoJ2AeeuY0I/
IUa7qOGSyCSV9HtrPjoH+sOYCZpCZ6P1sfDSAvWXmMVsXC9k2Ar6NhiNrxjQtn1KLEt0+RyUp+E7
fMAikQG+AEJdh4zwDEcaG1M8BW3KcPclfBYkL8kxii0C3Gg+2UffBmdS1wN3W3hJZvqELnI/kUC4
RUfSApkZ87n2zJj8S7J2II6rARwX0Dj5f3FSY9mE/KxZeV8UDd0sZiS2/AXU7PNL2GzR0Bw06LTs
Vj2v2gqOvfJwfXt+mCfwkbDpKRy43iRVIDrDH+RcXrMnsUUHnU2Fp/FxsxUxL87AsTlgCOZ24trB
uZj2jjkJSnXPgnlkivCupMeTxx/LvfiVTVAWjL9Eu16JNMKVKiEP7bdke2TGyolUDTvZwrKA4G1u
JjCK08uu9Whs0ryBnj4E2yDOBqei64f0zjSr31jG0x90VkhxoGpgDqhWzSFb1lgBsII+7TX/rI6o
HkUI6sxalQF4PWUg+Ioy74nd2Ywp0m5xPfx6PWCVg/8mqOP2lI8bt24p+/dJ+jYz1Kflb4CpX0Cg
q2i2WTVXBaRI/c2Nk7DhvOW63eUQE4mXepNMVs/IvIUXNp28i2SD2xqInbYiku7RdIsyLKxk1jlj
kMzPLLeE7kVnjFBPyCYtOVH8Kw8MhWZQb74KGnMVvIP/YUDKL1mhmlJ+SQxrwbxkf0IVrMkTBUsG
X+AscOg9eJwlwv5ySGCgiZ8hrx8wlWMBlN/EnqJspVvdJALI/R2Gqo9kxbs9Y2JyGZVYHSECFaKr
lsfZtzSrsGR1zE3oTCiSlUuQaxwOee1KYowDLLnIoCtE/98yfjbngpSOex6E3eAAZMfGZ9ynywJo
+0LuPQREtSfV4NhOLqnE49bw8tymGvIRKd1zy1tx7gJe2IDTjJ1xWTAfiyzl6QD6Nc1En9zpGfwr
h10wkw017+Mza/0qbzdgZNp6Nfdl3alf0OlEmmR0dRQujAo8pXxY2mpFrtpHEu61/eaZap3I9RXF
dHKtTpGHGBOfeCn7IF+RH6wG/pk9+dLdF6PgRjg18Qasqf6lttkz2gPW069Uajii6Z7/u6Tr3xGw
BfiDXINSPqQjtGZ9uuzYj0dA26KX15cSNp2HkWBJmY7fH6DQrvT6j6O18HYgpYGbQnGsgXygTnmh
ZVWh7K0oP6clQnZ7IqXfVD9dfKe22piGNJsxuYDHJn/UZl9NsD5ptlRTkOBZ0zccQY6Ho8uQ82eS
tSWFY/xPD+fkqdgse/DfFERabtrK4XnqEZZK6dFYdIFe+i/3l0yEhJri3d3K43sbppUGuOONEaCa
dynkIHM+a6liy9jZRk11YL194Kjua3sOwiVDDphuT7C1G9JFl8m/XIbzVUYImqKlU+16o5bsareH
s1P/9rHcmIT5DX6Zlxxi5QSlsnb0YID/TyQrMgCNwXXu2IAj+YnZdMdG9W9E8rZCZhPC+FqVZajc
/937lTZH6OC/o6lgCM8aHr9VcK/hEz2a32+pQ2S2DAuXubs3sE0uUC2PtD/RaeRvspxHW1cHWEFJ
jatMUceDc2m6ePNu07Yym5ofsarEITueKvZHknomLVDpHAJkTdAXfvz+ew8foHZitckgXjfeMA1/
U+0qUoJxcRu86O5YJBkA8LTTpRRfSt1K7wi3hYPzXzvbRBSuxBP65txgfK6tyiu+EcpWpNCr7GsF
0l0VzfppBX9JnGWfwRRlAvcHIVOYVn6ZALfxgbgG5xETtgzS/ehD1jttg+WNG+P4f1v5cJtJnKSl
/IVYO/K2uSgfgeD7mKQ2X8NkcRKJjZP9JE8bU7/u8PoMiPFBqZbHOug3oLaEyfmsXU4zMVIeYtFj
haZxobaqtNfjaIalZkPdqmzaNycOqHCyRDMtMqSvV8r5YjuMb02jSMBvDMnHVPuCDcYo0L72rdLy
Aal5luYRGzVdWGGWkmcsiFXfH4lr4pJxi10APRgrCCsAoEIGHPot28uUHLGPE4FnqXS3C99uD2xL
m1Fjp6VXTdbqq+tDLmqblG8JCpfZyHiiah8pAf3TgVo22J8pEPhiwl2KyvWRA2sQlR4qRSvp+8uA
YYSaUGk+sgJGilO/Pn4h3oxKfMCYjtYclo7Yu+9P1WXfFFb59fP+ULKkVCE0wp30E/O8/WpliB+d
cfbK5vLsnRNhtkCoWDoFaTTBvaCO5Nnxb7CN4s1PHBvWUg0WSl/ZviiI6kYvIDIwNGPre14nOoLl
Mj72Aj9fx965wLnQHflAi5LkN0sn7XvJfTDk1jByCnUJSwmGWRl4/RbOMIvc/2bYPbp8GKmAXEpl
IaeEDHD1Tb5gHGIEPOMFnFq5t64tF0YxYUgn79GNye0JeuTHoaWWmB5Vsz+Qk7Kr9UP2c1u66A1y
uhk8DTuiS9b7UJ+QcGBCV+Rzi0bM+ivuyCq5yd8CtbknXc7jwKQ0cx34iDj1j1P+O9nTU4tCQ1VG
RuD/jnbdKJNU3MH693iDrUNXhS223SHuB7USd1Sgv+ZXLyZ2a48BYsihUsjVZsS+8HwYzigyCoVK
h5bXlk3iuj27xUwxfnOilz0qDWcSREu4kfwv0MAHh8UQ7lrdV00s/rjhD6BUIHGWH7p/LphvrxLu
48pJ102BXiSBDuTKYhxPce+tX7wt3WHpO/tsbahHz0AkKbpGOFPgwQWa6VuamXpPcUL7xKN70mEt
YeZxEyelB+veeWKJZOWjIGAmfWutTZQI2SVyU+kqpDKIShyberDfzh4QPoxxUyKLJhr8ZHpjm2vE
E5olrElVBy51bfS3wuHEfsP528DYVZdRnz/4m+QAvuc1/KBEnhaRwqsi7wrJSnpSyE2O5mfgClXm
kvzg4OEn5X/H1Vv5aha9TqQc376aF9ocEqz+XJ/vkaZF7l/5NQVVChn4Oymg1Fn7HU5s7IR7Wwhn
4ndFpbLIzfryR2RVUh8RffK6Fb1l6gbbfghRbFILa/HQ9xI0ePWS6yGU3MeJOsFGB9bexzFzNcFS
WpjsNT9RiyccFMbnf0qEqk9Yo8Oq0NgkiJ9ZYmpH1+utAg4Ab3QtDwH0YWLHSs1ZyOy/7qVHoEZ9
DgA9YyrGQlTRqBb+0NeArHDz9AZwQZHfpwcrXlCf865XN5C1kz3ihpjbwVQ2WKLybkC5fmLqJp0O
iC/i17PBlOlk+eXSsL37TJ7KUGXkVYlBEZnQpjoeGMSJsD01JFMmGE2LcEnLRnxmDt5boezOGNWe
0nHjReNvs5v3/yWdsQR6ilY0PcnMGpZ9UTtJcbUwTsOYKmZbVT4gdl1UOPCiKjg5IZKsHKIz0JLJ
EqQIK6o2tYv7aTM4qakHLi82n3L14n4dmB2gcaFlv1kqJwe359r2M4FzDBX4WRqQxUi0jtVzXhsQ
pr2xetyaufeo6wM9FKZ7IlujFHqIxbiqAoD+iGRd+85yGpgSgQ7ONzik8nO9om/2jF4z66/DHBV1
+dUOvAthwShWP2aBWWDCzUW/EJcHsTpz4cjALvsooynOLmlrRGieQDQej90RQPJM0dmhjDSZJQD9
E5mxALkFUoe4ceq63XUfyoD/nFQRBXdq70HNQqiW4uxIdngx0VDuFe+YScvncOTNjk8k+wZNTFZk
yw2gCc0xJHCSXXFGYv+ZSwOBbsnTnLOmtlBfVxxqStDVetEpAo7YOl33GhWtE4hKqyVYh1O+Cq1s
GvbUsthJZu+PUjD+hWD15aKeWOZAFjZVfX6RLyRdy/lmc971CIzRitvv2RQMKeM0VYbWEILtZZSY
C18vygi7VqwILgrrXKm4eZZt7f5an77hGrHduOtThnsYGARp4WRJlWbWqDvO5FkSH8xTF3pyujLi
uzP9XwESHB3BfnHL9xmIEsrh/8RIkGjm8cmOvZcmzTxwdX4uVDXz/G0tfM3u5Wohstu1VK4JEe5l
mM4WWPFxI36hLt1qPLew3Criij6Ag2OW6dM8z05n+Dn5EKszvUKhRE5qPeY9cGlxyCw05jLnjRj6
YgYoMYEoXg73KVRxLhSz1Oy/NrlrOSI+g8WC/7EhIw1el7gEzqMI8aVTBzHzkZBMnd0a8MBYM6Be
zpuH32eeuxrefWcfxcnwEJZOzMn/Z04B+nkMpxFPnfIKQA2FqFC4XT2VtiuHdqEEKk8pj5geKpXw
RzmOFQolaZjAQ/kHTb4spjJcWn/c3ZFnPVucOXbp/Jvf09ya+KfXc1X6r2xrrFjZlDH85iAJcVXp
o70WNvycrptzfoAVjm98OkBZ09nQm8QbHIRFlhM5Plmdv6fWp6g4sQA4XmeNX4/b3qRqwOQbZ274
sEnNkrQ+/eo0VENAJRs8pjwNYvKodYhDTwL2GGSi52MuYmMi9zWIPLwhkIsipIF7o1fEn3/EwvLA
AGYXppwAYemXKr7tkrM+xQF+eD7bv6K7PhE3FYCrzJGFhCfTPAu0cwmf521iGB5CJ1Od/FDQCWoi
pie7GCSZlmoYJ/sSH+lt1KG7eb5mnd/0y7DZerGy6go3O6sB3owFbsyy4lYBPLEA3IbeTTLKZt0M
xfgig+wrIhAYouJsEq1nEixWloOkdpWP5xuqnssH+kE2Fevr0DLagK4LwwM4bThN5ou3n4r2X7Ry
IqtTSsb3fruKbaGuzX/HRsgRxmyPG/KDJ65tcZXcjE2LxB8ALQ3K7VCO5nKk4P7pPWxaeA53D5Wu
v54J3BUYtUW2oLxSRMrj5+QTHKXs/H1+pOIynC0smh6XIIwzqV19HGtbVM8AmKGNEWHyVpbhQUax
2ih6R3drQ1CVockFSfFpezbxuRAM0hyOlQNgS3zb+52IuiaRHlFL43kvZrKY1GhItWSpxsMkdFTy
DDGceJpxegcw2QOeil9158mKo9gPM3jEYRBjEc6ey1VtqVkTiSS3PbtFoJ733Gnc98T0hMIVGyBy
yGUOPRHxe42bw48uM53BEHtwAJtxzsmYb9eb17O+QysiMp782nBgOidDB0ZXcBqB+ep9rQzmxzah
OwwpRdRY9v8jrDl/t6fuLEFcrfjs/JPM1OYl2oP4yX2ArRVBIP06k7rHBSfC8Rvs2xK300I3uW2B
bGkojLNrI5kyqXokIv4i9j/eAZ0Gp+qmLxl7AciYcafA04dCUkwcNOlYZWMmyu+bgux/qv3eVE5/
DmQC4YrYXc6SDTmHV5hEw/Lj/R5XoFkNxjhT5YGzmKwA7lQXz7f3ac8rpXQ/RnaJ5s3SV/N5+Svj
6Ul7MZ13IAQoHXEIh8Q/DmkeNpn5MwrAqoKnZa1usjTGTqvh7lebHmF3K+LpQm2Gu01xcsuYLE9N
840ElSI5XphM/pMb+J+eUREbyhg5GGDlbzzEdgkq6DwhoZkVA4mqnioC6lVVeM8wjP4ixYqX/kWl
EuPrv9I9BeEuPIUUs4Hdl7BfCt8Y2lP0MgeXbBIpPkH/D9F/ba8eqI8HeZRe+DFi+dsI7t1fIyWQ
O3s1uhfUz5NHSoxEN+Nw5tAJbQGqkuqxhJ9qt3XAA/u1QDiT67mOWUVLtTIsmzEurEV0MFjhlf0R
83OkUOTj6iAPSWhdChkaoK8eD652ZSphj7N6F+mXrvQ3/0oa77wRYfgkhmsMPSq9qcnRbgTzX7mM
xFaQ9XT4Re4Xl8AgVQx008gToTIQSPM9E3TLqJIAJEG/eXo8Mzix0yCXdsNPWSR16oNRe+QP6Hms
VlGo+DzQAzwuPez+gwFVxbO71mmz8Wj2VzFthJRhQYu6LxqbqQx/SVr6HBiJBHfnj1Lhwuq8ywtF
37plPIXr1RnSWOCjAe86hxo1HEZuUxlpyrCEeezjIxA3cvOaInuFuylcPT4HS0tgXShtxnWshyci
S1vc31TQi+MCof6/eXDAQ95XKhjIdCIZeeB7ijH/dEwk+6pekaNeGU71E4vf/sS/2ltYQV/MZDc9
CQeHj3q+4I7AUK/T5uljiGJYGCptXBiaMdsGIfhukynr/CvxzI8z1GA+omKodWtplJ3o3x9lPTVc
LiZOMfSDT5pXAjXDm/cxsiyEZEWsXlVyGrFZ0YWvrgRs9h5vRYtPDHDgrpZ1f1+F19+dxzMTnXXH
wfEhNDlSskY/sQH5+pCuazCAeiWaEh95saC9KOgEyHi1MVqvIhME/uB1qczgqOOKgw3cliB7pzKm
xoXVXkfyPwCpS1HD8n0YkVjk11sj42eGLnTJ0IhK7FVq2J9B2V69knedB3tius9TW0sxjMfQOX/t
ln0t8jblfhlVSLg+OVwDexU/f9pPh/J232Yuar0DyJPeGogmC00/sNzyD105QvDjA+Zma8+uMEzg
RRt2bcVqE0d/1rMSBG+9VeR5gaK9xqQrE9cqsu4QXCFDuPZw87/yLImSFkB5adZIDAJg+QbclYx1
lmvqs7LJ/hEINir3WTM6RPZ7n1n1n/LejuDUe5TkPGcry+bx+VrmUYV/GL0YFZKRxxtA/w0TT3Yc
ZnvBRdqnHtretzdtugQ3XtqR4L0efVhLabs0aiFp1rN3cBFo8+uTq12XVru1347S6AO4oFaJVkCp
H1+G1SnqxxWm08akiN9t9Lo1ERaAvCuyBkZoHjiWFL5Cs9Iw+rqnQRt8g4JxPaDR17L9Kx7jlhMt
dHOti627RSstSYVS5hgSQM/U80P2h8hbTZkoheSMyy/gpf0g+VYCmql23zgeUY+ZuyYN2S+LKtNF
64rdpTaecWUkwNcHHJlmkhmoGgaMT9Wf6uOqH7jXIxvidAjDsrHtlmyLkhqswT1St+Wi6+2C9Zlx
DHU1ritJcP2iuBwEylrHuGqccgGTyJkox5b/7borMv0ziqz7+1aAMYxdzQ7N42Yflwqqnc2RqwyX
NolJTfPwyUDs+qcYIQyR6l9zUSz36Fay4UGbtOf8Jzn9DZ0EfAc/miovNw8HufF1o8oFBBHhZkg1
ejaiK+MZPXoS+UFbq6SmUq3j9zH2yc7Y26wLn5W8U8inVl5lSJr9jy3Rqj5EdrgwiZ8nFsfacYUR
cCEAn0q7uZblljaAQQeKbMscoY20GWTRVAqdNV3AbunXRWPbL26HiFsg42jCKz8sjwe0YHIBxeJu
AsJQcwufIoAbS89h9i+q+6F+KOHB7msfxF/Gc7QwYQ9DLL0NQ0UiDTOxmDZrD6YS66zqOCbFSAzT
581e4AvaL5MIaVoJazwzyWOcf/EQhLmCw/Sh5BLOKuKdckOgQ4b7Gz2F3X5QvMP2yPeNAS2qhLc7
tBL4NXZe26ZW4MA7f1hfR6TKCpESIki4ehb6uNpD7TZ1AxeXlDupZX8thpWa4uTPWrmq28yWCHDE
tPoEcDd2XNLT0pPR/6HUACOvaZRWRJI6mFGyVSnjTJFSMHCQ5Q533q1ERhhHLObCRIPYpziepqHY
WMf4tEPP1mG2TucIiEcxShHt9hDurRxJm7AryMwF0gDGzE6Rd6CUj0e9qmlPCem5mQODzUUc6vEv
dBFtVSRTXORb9e1cE2cTLXqzoQQk5r2LnhJ9Bnm01AVGfQ/OSxs0drvgYnuadClZpCs8WUGSMHCd
xur5cBfFlHQxAchmfUW02UoLOUiOIt7dQ2zbJotGEZxwpNvcGMj6or/bkZN77FsTyO26wY4n9paZ
b7jqMJpPSHrHcytdbkuBzA+q1DdVidNuSRwvkaMI+5wt7aXsJom1d7Ou2ni0aZC3APhYRk7P+6XS
b9Mp+uAY/+rGCVzMbWP+aQ8bN0cyAZ19RqoVKadd2/h6fxL5xu9oomEfStxjYaXppYgqu7PEUlPx
JOv9MWU56dwirqz+KfHM5pMewHGSHWV+2AGI8CajvdswDBWp376QaSTnW7u2YrmCpQCUI79fxLT8
s7GrNMX0xZphwc08lfx/nWwNllMKQ/KMjXNgQeVC6SxrfMEMCvjEfsHnyDNXbqnsayEdSZdHuMOK
iNMBfTfiZr7lxmBSEDN2K0I9+Xphu+JVNSbYs27iGsJjsfxyrioAcpc7eYK/Gat0dUNYvLtEZwEM
qDulGjNZL32uw2vRGTEOKgYD9LHAWhok26JGcfLhsPYVTty9MjJ/QZfSams4ndzKpFI8VmbPu14M
HD5nJP5yNNtC2iuXZgfshOfqmBztrhyRzSfKuetJ8XS2pBL8NFQO2X7/LvRIdKNSrC95Nw7B3juz
aqhpv0uAcqiUIqc/tuYFT8WOT2k3mz2vmPLXeBt5RefgsXwro2FkOEfHsvg++64ZqDrdAfWUbh5w
gQIKEX/n6pZLk1r/W6WH/K2NzWnu0MSye7+AhN6yXHBC+zBjruVfh1BM6tbECOaC2t875e5WNMVY
peI1YlJUF+ViDghdwrW+/Eg1H6aDsjP7mT7xoZ7VI2FzubynUmAd71+OM03r4AVWTQ032R5O6R6E
iNTt1pKLcCa0S7PMIgDJljeXGGs5cj4fE01yh1UjDl58fjN2w2whLSoglzGnlyjA4L7IcKGRR5Wi
dpk4MIl0NxxgHWl7e3mvlFGpCUk7X0odqEanq0k8UQBUKkHEUHu1G91qYXcnvsQsFDljrLqvZDku
Pz1Cx8kXQR3N7Tn8gTbu8KeoKMHttGqgjRKEMg4Xz4JyRSt8cnGwb/L/Vrv6UztVd92C34a8fmy6
FplTDqYZ+9ST5+KiOyn3SewF0mQg3TFE8s9o5velZHSwMLeLs5raR0SZ5c2AW24hkLuoRvYrzIM3
kTKlvVTTZpmh0bmWIxeitMwvA88y5qsT+W0v+7fnCDsGpjQ81Cns2VFsedAAa/Cq0FT2f6BQt92n
AcSSRKoWC6fV0vygZVRsyrBRD8zzxDc0rB9tl65fGlPQu+EeQ81CFnhGXxHldavRqkHvB/SkJDCX
IzlIjNKKh79+xlM2VFzZUbcjgCN30eHakRghw8X3RrS9q/D/aAJ+wdQwnS5GcNWkM/lgBYGxH6G7
EfCcGXuzzgjrMk/2GsRVzrDk00Q9PoeM2RKqjT83GbLq3yTyzoJbfjodSL0dSRR1UYQeBAqlyXEn
Yi/7buHVk24rodiaxyP/llR0M+0LOlwJiPvicE8qaQFB4XJL6FmfJjvMu70o92F55eZnOTS/2TZU
7sJ7sLOzCCVcdwes3sAeOp9h5qrLNbhlIbz5Ohh6BCcu5o+9vugVTVovqJGiEUF9wQ9X1nFFEJdn
xd2xKBMy9/vkzgut5+cWXtu2H4DxJdh+qImrl+932y04TsnLLymfrQOfHwK2x+zf7YVmZS9xMxOo
kEhBImFf7Z7YJ+Y6+BalAnT93AIwa8um/X+6I+7rWyZV0Q2aVxm7luew9cznd261nA0EulkgTff+
p8TmFXlkogy/5xnV4iZHSPFcw7fATBD8JwyniDd/CciXB+wqwDUjrxi4aDh35pyTFaBsxmTQvHgZ
pLh0EWVLAaWSoX/lHzlEuzdqpoNy6rCZjCZhLJRWWgtG2qBnw9wJjHvYbgQEpbIT+ShAVgGDJ47e
/RBXPxiWzSpIHAe3zn90/k6+Q1uQ37qXC+vFcgvaqwuTRbPGqcInsCAOms66Kcadu7Mjb4zQhTSE
d7LwXcvYf+TwvM2PvQecIjpdsz3epN0RulOju93C571La/pb7T9PrJ+bRpHxgB+AlxkFPpmXs6ha
r231o4wFPid9yfjRKRk8Rqm0R2adoJGVGnaptK0oEX+47sN+d9EClcdcB5fzsspa8oq00iV2rVQ2
4eD8tyA6pXq34mpuu+iDgv8a9U4T+n79L8kVP2KG8kNXU160Gw5GOZ8n5/bNUxYgq0/aJNpMGo2S
SM3dYC2iHuDX2GOY5kvVzYd7l/o52Eg9MiC2Dqc2xux6AynbG+4fed90O5wNkHri1e3lHzlPh+tI
30pSgOsgOR6awiSDWH64Fb5LlAGXNXmMLf9nBseVpO/j8A1AidteVXuxwwbIMkjt393XrklA5aKw
uarEYogD+MjsmmEP1RR5Osys8832rWBK135gtHEqmHUiBPA9tXxrD3aD9xVIwTx1NqDSLQyjbERc
RgL0KQiTph6gB2ZSAi3Y613XF8dexvQU1RMnrUx5BYXelFP1tH7ikn3zzfKdw5qlsHYTQ8QnQgBh
J8lvn5oKuZfDlkMlh+u2YFDimvDcmMlrLxcc5H3c53QjxRveqembvJape5jRnf50XdJ4LYVkZjyK
AxaAbeJD40uLJUhYOu5VNv5cN6GGM7cSzFJVCu/s9pV7FuS8ygM/PyOSTN0A1lpcTS3prgJ2tEo7
XXfRs5J7ehR/Fi+Pc/qVUtloKc+I2CjmgOwNw1USEEcwwaiYUpajGqTBCxmdmteAy5btbsNY+ueS
gA9Z9eAty1EPTqbmk0XeS+c+wu0XiStr7I6mVlIBy2mdC7drbzHOoYx+8ycdG05lRRelHCHlnSgq
ijGvB0nmfdyUJdpifA7HKP1ao+YUUgMyNC+VZRCTC8bPJo/vPPLu+mTCyuBl37mACIPzrMNcx5w+
LlYziwH5VS1n5enmss/tDc/dDLWmqugvAg+iMMJw0z+iTKPkUbf5z/KR+tmMdftYG8Xf35yepo3w
grcBceEhbkWUGxuJt6FZqjyTDnz3opQFoCuGuGFkWvTrdO56alsOaFCwX7wyszt58qAwbZXp6KX4
Ygq3Q274vFCbRxjf5vGDYxU3ABAvdOtzFxA5m/NQB6u+E6XASQV0hmY/Gl4o/NuQRCdkSwO6AMTV
LwnQr2wH8d1IJoSvVusvFAesET0BtTwy5Q4Q6dmEt5g43H8o4YPgKZCNZtlPyuKidd9Ni5fprifJ
NSGMmMCg3J76Kyxzfroebitcilmp3k0Ck9M7m2ln+Y73qqNXWdVGgnGwrOTZJdxKY/BLEUcCieYQ
dyrKIHSBxe/3uXiZpGJtA0PO9M0W3u2rBPSiMLSLsyfjae5fLzL+ggClwpv4ZbNW5JAYt83/iJW7
ZnMqsyPcBfZgWQJxLpLuEAfBIdebqJlBzlT2qyq+WbPX71N31ej81zEITnLWVWijEJ6Vye+RzT9c
fJFUUJYR73v4QjuGqjqfCLtENJDayvZJlZ+dTE8ZkgTuK1ix3TRzvbtCJMBKOwadegZ/71mGNVFU
srF1QfztJ3ok/4fh8fsPU1QZb5Nym2q+vMWr86CI7CRew1Sa0b8QLuoSUsOpB1uSAU1Dflwvh+Xw
cVOuRhLODg103Eb4qT4Gqv0/spNStSFr7ghNmFgj3g1nxMrt7cVVUqKo4fzUTqWdNjtU55eVtoMi
tz20YPnIaayD2139vYffGCeurajWOOisoCCSfGmUqs993ebMBOaK6WLowD/ycU+oBLCRIBHA9Mu1
+CHvRCQvsZMV1csoL4Vu8fvL1Jzml2eAhed5M/Gi9o3VOd7rb6W4sLXO0Bl6XSJduQT8PgEaNBpT
y6n8yyXk+MVt6z86Ex6H9jXKtyBQoH5a6m+TMo3BHKlgUQffYN7a/RxLMCZ6nyVlwyRabgkuYYUF
MCXzuNiXVaLY8Ukn/PN1FtcXNzeSQkfpOGF4Po1G+WjMDj8TBW8PqnCMEj856QXLSE3925m7rCDu
Iuqd91hHoXwBmqhJPFQdn4IGYPI+uoK2WUgCnfJoObpJgfTWlY0HlrIk0zvR8syj6SXDITRIT8W5
DJm/RVUIzX+Y4YVN+VKJynPNBxeaRyQ0i9svzQSy8+STqsOijab6XpBq+pT1IgIURnLI4RZq16c9
W4IxE+kbzHwa0OPQbzQ7mPjlPPo/CfxtfTLiti24nwVJ+sOwyPtQaxopQ4TGy47XGFFxA63bO5Rr
FUb7y+dWC+0lQjv2db98pk2AgwgXCB4mltY+/PoLdOW0kuNrvU09n2glPdAhu5prL9RQYlC+v2MO
0n0Th4KWSb4McwxXLYSSRa8/cSYDiASoDp8s+H9UBFasRpS7MjsU0/H7QaBgp6X7rtSQhpSSkNS5
YB+kRCQtMTR5QqSZ/rKVPnxPA9lxUgK3xHP+DM7UQV2xfA9yYV56dazKW+bt6Qxqu5Ie4zQZMz+R
ZlzJxlPYoKAFlL0ja7Wp23ZqG76vhdV2bYrkvfthoQkTNb8GuiFiAJjd5fwoKSpBzul37jjB5F5n
IsQDB08A8k8X/Tf6hJwCJxHuAIeCWSQ9cNzO63JkDBJwCIS2m/gVKPIUymubsKxqcO9pCsEWS/Hc
j0YFNnG4wnfFHiZh1jVYyITme+ttAlVQEf3m3XfD8KL6Gw1+tDGJvm2Fse4l9OEcIW1uGQiOB5+W
pNrYxBVairBuZsY3+Ead6yb+8h6Zy5Ix+Ix0mA4O/B33TRhx+OTQLrX6zLJ5xqcl9aWTrQpxTXYB
FSTC4Dc00RWNLdCf94eg3807NQ/N7cUn0iZ2io6JiYm7aFcjBGnd/zqtxhYPLlyNsG8vAt2a0ZTS
oi8s3iGAGKySen7CCZ19pElbiYA16lenGDPZTRXSaGurmoktZfInEQ5rEjIusyhrWglU9xN8G6Gl
6/iD8rZFDqRNqSJcAYBPjhDULGKPlBIPIMztiN9TWSlKI0KckJJUHtZybAUnObKx4GiAfVy2qQL7
tecQGSmKEle8rOPUeIE5A3rRaoqcOvJ1EI8mzdIsLrEV081m+t3WVcWTlPrpc8kMNmsGmVV5Rfdv
r572cbvW+hLPLKbb8hFodLFpLeEw/4HGsBeSGnTK3JwN6DW4Q+Fd4d6KFvvlhZrnwF+z2zm8qVxN
IR3+/VA2zWnFh3DLjPB1iv7FRLPHWH7E+LfRyjvVZv9s9vEL5KNmuFf1AvIlWW/qPQnnVQ4mZq5Y
iVMAkrquYhE2GsZnExKm2+RuqiWNzjkhm57RrOIDwQ9f43zqtF2BgJ8vRHkf/+5fd5fsg5l8KfVn
bf90pROrJm2QByolpUZtx3Oz3RJhDuN8QZzY8X3mkTu1hjTHVF+zax73zBMNq5SX1rDiXvkzZG3k
XjWK+dKC+UoWC5zk9TcgCKprXQDitYy+HqMgsy2P5SevQJVuEz3xXR+k5BvvBVKbkxbiErb9kXJj
B3bue+Xsmz5sgYq1rOPkK3y0hl9W1BT8VVcgs1bX9jaO7qUZlgHj29ghn0TUK+zbpAl4iqAbSeF0
07kRKvL9QBO4B0R1ahsjevh39A6kxoNy8xVYIShawalH5yeXJrcDh4NCiV5tXXGA2uxEfv2tU+1s
7qpATQRxWmWT1DkWKqkQ0L844CfDYa1GuOyFzkPEcf5fiDQCswX1R67Hy7TNKXJaYNzqia3iONMh
Hb6yBg1PDz9g8LEwPRkHHI+drb1vU3L//DYwG7tAEFSLtlcLbwMsLSTeOAlAn7RGBWvr0LZe+Rtg
oxfCE9OaDlka1aDfv90P4HxgQ14Xr4VlPTJxaGGHcrrIXw5KP1NB8tozlx1mynl5Iz2guocLVLFf
pHlJYVDtk/7hSPs8if7t4JyvBiuhDf67vvF3bu5MFVU0+ctA9F7njvfNPra3zxNnXo/7sLGLa3fm
mVQ8CjrF6Z2Km8wBqEhOEvhS/Tmex8L6slzKAovjwiYyOyznBuezRKVV5MK/XwcJGHLCFFKKfBlV
o5IMCEo7017lLmnpr5TSkoHw5u5tzZEzYFwGC0TiQroQFa+aZVAt2tPO3ih+K3Sa/prsQaKecogY
FrykcMTDr8MKfW8rCt8wgmnPDu1Gc79xaU4MdCH2ugWJAhi5TcvaZA9E/ntiCVjkYc/WC2bGgDcF
Ewe5Ppma7IAguOLGl3Nc6G9LbhK4HPT2DVawKHgkMvCmx4lwQbQSftx4AemY5c2fgpeNvVcOYxdJ
YK3ysFu4qpNtJr63b7hoVMd4TVPgzgxQ2cF+rT48Er6imWc0Rqu9+KvyTYDBse1Q8Fa9RpnircXZ
sVh6NPxVKxyvGxSXjMq4HgmqnjSEePSAWcfFo8/JBV50HfVcE4nf8CbLmFUupgbrxCdqieM2aWOL
oqSJf5Zv80H/YAoksrm0nMSjGZe22t0VDKW7xwHL2FUZdc/Pzq1uL/jhnNr4DOXBv5m0Nbgsfx59
A0ll1kf87PVVhXPdmvzQXogLb6Gmq3WgfOmLjOE3L9RiAYJWxGsdwCGMuac4ezUwlJvJp9RKfeNO
e7jEJhmqtDYaIfxPJH7YTWFwHXBXl2xY7yNCPb59t5LkVyCOusBx5Y2Dna6jpd1FN4cG95lJjsux
UpUHT1WcNyIYmTNvh+UwCsGtyLbD9ubTZIkHO5Hsq9Q2NjKWSEbZveapV+NwV+hgBgWNTxOT3ECL
Aa+fgZhqupAJnWsUGB7Gf9MuI2IqKrtOppO9Q65ijf4qMxt+zGOxDK2xmU8FY/DEg0MxZBFWtLZu
N8/i8euE4LCVDGBDzADv2Fr3GUjsSlgm9talvoo9PccAQbmAVggRBrsreHunaptdazBeiTxEqI73
EfC8/UrNpIBGVxOc02vhdd6Vr8wNYl4IlMwmjM8PdyoBVyBuCmsgtcfirIFtSK5yJxHLiVldqdKN
yqngchmtXqSsJzqDoGwTiEvaLXfo/3Eesp5/hmAqjbVaI2Hwg1tNMV96ghKGwyoxpf0UTClAggcI
xZYnWy311XDxdr6+vS2gnmKz797ApJ0X3CqiIvVtxDmZ532II+CzCUpUr1ap+TwK70kPHNMifdzN
uewWa9lxf03EaYogCbd7KSdQ8LwMJWbhJsws4WdJFU/b4D4ynhAS1Tf6p/6OTh7E8Lr+JDYKLD5r
JBTc95qSqV9nv+X/HcoFOzVtE/CJ614k/J8AcwiApLzQJTYxVmYaolJhmHgu/ljuOtC+U/mTFIKg
TtARu5DfY7A/SkgoKgHCtNKN6Kg1/VkQvHzAKQThH93ElyEzIVwRYR14QMUcMj9LL/Asm6XJUPbE
kdC1Aqz/LYUkZ/x7o8Zo7R7WWokrVAQxJrAE/afFuQlxAEqdc/wzZxnnsVTCk/MzGXEyl9MD5s9R
bGwYY1M62oAy9Ovx1ykhB9w9pIOIFRJBh0Z386kxG1AkUtsArUrAc+Ad9CaS7RFXPvO5mF/ldgkC
uudv5dnP0o3CvUp3LVBYYYlrb8m0ti1t/wiMcZ1kpNEg6s+eSUNaaU4ff7pLIqSSzHAJdGBQ9K2p
2BdxH50oT/eg4BOddsO0uMmjZeLJgbF7+6ScR4DAtPJfzxJE+6RAfahhhSZ0MjVmMr620fOkBt1w
Ph7N4rFoa8M2yKRDyWi2w9oNFb+96F8nxtzkng777lDnqqaF7KxDVGcDlHDHgvFJzsaJH4pQ7BcP
ovAVM8xPzKQP2hYuQa/qzWhdJWX4vWY/D8aBhccWv5aDXjKGoRBPUQDmPqrvQMchuFnLO1I3GYoY
YGHIMAVScVyST9c7KcmO+LHlBxDG4V+gcgF7lPQ69N8MbDowQLAwL8Bdzoj84kpmiOQeCnrAjrv0
CtBCEMiMLtuBObh3OQNZjkpIcpvtW5EuWTtgiG02bbtv85zv4iN6gB+qaOuz+KT2vdJo+TMLgUdR
jpLbugenvpL0oma2wuvhKdlLYjY3cwPhlruEOipIKlQZV7H4F8dyHq5lInG1k+CTZXA1JiqLFEeU
qcmfa4zXqgzw5I2AyGizofgVoHOOrz80CsyISLrB3/IS4S+0roURZtOIgcRH/bkOod4m2eprQ316
jPLolHOIpTGtGtr5DSTT36btFI1GibtIAfFm3i5P7fabkDLmq069BKU/qZ/lv94luTP1Dulxn710
a40HX+Wdl6Q7ozpr43Es44rraBB4RoT2QYZCzlZWBf0Cd8bI5ODwqVDjmEU6AFmK9KBTZTRatTTH
HqH4dYZLjcwXsmBG7eONv0XgJ9LknwTt+eLsaqRD2qVl1f432typp+7AlMrAGSNsQ+vCD9hM4mhm
pejm5Kiryk5yxdLL3wJs6KHSO5ljgTp0KQMrncCk8RDzL7ewnSmXM2d0RRqqtvYMkvodSrWrT5wo
nAw4C3iUyOBGT7H8S5W2XAmFM8xQ9+c53/EC5vFvg6mCeKmBer306kL28o3BU2kCxo6wXr4StIVX
lrQJsL9QhJrNMU+7YKKvgP84QAc/x3XOaSjWenyiCEexVPwHOpop0Rgk39Z/ByBBg6XshmtySF5N
vNXeyzzTMIszcB9H4fEODLLsv1EzRJ+F3FItrVob1FRb3f3JBQMigsqrfPO0JusfbZOYb3wilAjG
S90Ch1qqMJFO7VGPDWI3ruX1eD08UGWRV3x3wm7dVwoFEIz/f9YOlXp7S8SDPPKEXPbIwI4RrlU6
61hqenjITlVzNQBoamAyC2aPQZkB3hiEceJe8f0YoUDqObUY+Ec44fR2FNzsIcOJzqZJ6+IB6r9u
GtxBY61iL6/3vCI739wFPq9/ehsNKk/WNivfajwlPQnK4MddAoeQ8ynC+nuvcQG+ot5j7sZw58QP
/IQoFqNxxy/ezSZzpnEQfbatRMReRq7uxQk31P5ehaGMQmiQz3DPxNGF9U1VJk9m+DAAuuvln/oZ
Rrf3s85Qnm2jMHe525OLPB1mkqmVbsrAtbUjmZhDYwQPd4EiO4DX/Kcgd+E7icjMGjoxNT1qYVmL
qnjWLy9bvV8AboG5xS3qwt30YqTitAZh5QdPXdIyJEtHQ6CATLtjYdYRmJCg7vf3/ZUt4C3g1/Ls
0XYVjH8V6yIX6EMT3fQ+nu2oEs1nUmzE/tMALR01A+/h69XAwahcQxuPlTYSyNcDNE29TRmD/bqN
UvendCljnDAcYBvmi6lFqSQyU11M4yma42aafy3KKnjqSa+SFEf0h0EHx1oD9u8K/19X5vATnGBg
+/kSvb9Gy43uNyfcnD1oL76HKI/rR95XvJusy7dFqo1BfIRYbIosFyIbhP0rU0VrazVZrkdvTZpj
yOhBEr5UCOU/BYhQYcLN9IbS+9AT/ZkOYtEspFFNiIBIu96/QPEgK42U3diW/3FU/fIzx05M1Lkz
uqgVXoYsjp5CFuXaZqq77xgB1lfQAdZu0bocXkzh281C9F8PYR7FvEx3rJiyhlX4oEoYWVDCt8+v
cvavCwgE3O2SB207vCLkdAVn+RRt+CgK80vuPludsYZ6VdzWGXWkvnW08KpZ7uxFtTv40YIw2w77
tBjkXQhUrPMjjWhKxi+aQC4emdEA/lx7qYu6BWst2+Pi+YIUvQSh7Uu4eZIwFJoAHAlmfRhZl9tv
nI4ShkpeaFZTtwL+071FCHwc/mUU8aPwDwy710YnkW+T7hR6KQ4048QfCwaUHJZq668Z62gjhPpg
1ql5Ca2WJS8nPN6aiDAQuaK85nO6texS0LqLdcsJa27hf88q6pQVMzmBRNCO0441Mh8fUxb1tPP5
fLoftB6VidtJjMXOLh4Z7udWrdlA4gA1tWx2BcFqoF6T9Sg0iUhz4EMSPVafjZsfv0T8KBz8yTAj
U7bYLLVaOVILpcyYTWEI1jqJbAynXZpGhoBCX62N5JiK2Rue7BZu5JDD0Wy08l5ElGAPQC8c8DyX
CGXHXHMtLRArNp17GN/U8oTaj67UFvUFYVctl1jXJswHNjwdcPEmg7mmk35hrl+vTbpUc+Mrzye/
nFeuDpNOx3wy6IeHKxsRutb/jBi7otWMEZWaWGq7Bji1ceDg5eMpDsxTKvJy/BOsKJ4idaOd/ZLr
k7vPTpb4xRvJJt6ENoH3hpNU+aBLzDrYCrnqj4IKlVcR4FvIh6iLBnJGT5tLVGllHIqWyFlvcoH+
wP5IZ9vhEoE3mrYNJKak+s1R/mR5ggSMNkWN6hghZlUJUGmBt8XAs2REy47DJd0GtiCmQg6XfyFu
N+itT5STOGmGiTJ25DhrhkUxiGkR+kd4PfoJbha2Utfb85bI8PtaH6oTgvX+ihDXPjsA2Cw65WfR
D0IusZSzWNEwLGyDxJM3j9EoYrp3LohnOfyIyuFhTXR7W2sYd4WzycOM0TaDbD1su6HLkpXclzyz
hdI76CUeRx5MND+UNZtJEtIpV2EPeuHujkN2rvMBm90pPoCprf5Xf6UtUfN3+ISTCmxYH+9GRm4/
B/C//DOPlJYKCve144Gka6jWsnD0MVrEK8/Svh6tc5KNTtKijMqJbTLef7UesFyfutV7d/qYALUV
6lAPlS1oYzPrM6/SWr6Ks+FkIeJYNIpm7VIWYQAJn0cgY85rJ4NQLfxltitfBIQxU7CS+gAH3EB6
7VsjeC7z9nk5pMaeg+ub343gjFLVBnbA4N74BlB9R/wufsgT9HSKXp2/K3dDcELTCrtKKRr+CFmD
XC2wg9zeK2YRPyP6ERvZQ9ZY99YR/NstzElu7vctLSxFbZkEJVD+nbUrXeIdAPYdBOzV/jaxtyRm
OJE/4B0b4554iJWm1bbx7xILBqiSkDSdGwd8CHWNKfbTjtvuUucHXAKEbqkKjs4VLG5Ghv0Y/whY
tkFRkoSe2nOLjBIqNVdVdy++KITNHgaeDK30/M2Gk2pAn2vGzp7es/V0JRDhj1wr0VjNQooCoXPv
0drDlcADXHtV+PzYoEfQNa0xH+v+gF+dpzJHpSr6tVop1Cg93U2q5kEFpIAj7HtEk9beqR+4s5gU
jw0t94F2d5VQtIOkMp0Uc1ESB+7qliNoRWiHpQgZZiNYzR7XHKLzf0ch+GHIzqw71za+PghHXcFr
+Hr4AZt9xYjcwM7Gb2o05MAnxsvUyf33gNZI6fjyty7C2/wGg6pbA1WWIWmozTsyyWyGYsPqVa9m
Nu2tK+I9dKHkxJaGIdaNxdOTy44bwHiop6JdhjcSshP3oav++KN7YOuRN765aTR3rSf5ZFClQUFD
AU8R0y74OXqaqQT4twHQhRnrV0+EbS5TlOlsAdLPMGvA6sdCBh9UqlNKDB+PFGRrCIxnN6Vuroei
FZMLpjJK/Jj0sgJJQzJ+cuB/HIMeMhLBbKTTxWI81et9hMCWmr4hA/8JA9VyM0lIzgiEonjBVVBy
KrtA0+BG6B282n4/K8XklJ5pNA5dU6I/bS/hwhm/Y6o1bOYrx4W0DsltxtfNb10Rq66OCVGWfQSI
egG5Iltz28xZMZ/hCrNEL+KlDD4I1RKFQaIBTCemAI2q9MEorp5Px6ZxCZbhHS0XFPVxsqiIKEAl
ZUv2+ywV4HycPh035rJ6nGZWPgBMwa/8cF2QS3vQKhaT0qTb7A70nn01ThmhrH/fD/YDSD6Q51Sy
07FxoLGrbMRZGDbNOEXaqjFUHr5moJKShMeWQjAYMxd5E8MIihlQzhzaLQLA3M1NYOP7pYquPorX
79qOhwESAY8ivJc5KTMEN215nCJRisA73n/mJ9+IaCCRNsVQPvKVQF1fqtz+xF5RrFQglDTRm/wF
5/Puog/Pv+mf+175NCdTL1Jcxe2E8yu9ko0sPIdVC9DfvyDIcJCg7k4xtkj+WE/PvBeJ8jA0JjIN
5Ru/Wu5hNDuDJqecSPqR3qe6xUNG8vh1QFS+Ay3P4NBerTU6MjW4KMsig5U2WdwauLmcDAzQ4AQA
E20B3yWcdK857Fl7YrMDZ679D42brWlGBMlUi7316fHMg7AcssqMTndbjfcibxbZmUBKVsqq853r
WKKRnOKgocfWtvbqv29XqPVlKI9OLO5OaAov3JmFGC9fEiBJxp9MqhEs1btebiwpq597Y0etBetg
Ojqp+Jue+uZKIyveWKvNkRU5upvCjaytfsDEmGd4BmJmvj+++5gbqcqUvMOked33YB/w0sNSXlrm
EwY03kPhM3KPIvyKaWSXcwMV1c06sNPkcDAbN0krrJMbqLlDCkYg6rZxAGCz6/Rz/lJ9ySI54pgR
93wxHrnkxsckkD7QHZB6Jzv19v+bzmTtDfW0+WJWn4FPIjMSrHfADJMjrG8kQ3HLVz/IyqIXZFwk
gyReShMf1g4DtFbP/h53SSreZR9hFCSl7hmfCtNVrf0BMz2G14VGvAnRNlNbPcyx2hJ5IDLL2Zdy
3/aR31uy5DktuAMPjeMIiZFyd0p/Wns1ErLwDkY2RX3xOsQfT5WJE+ybF9GqSdKBCH4yoc1/iRtl
vPSkdX32iXhXZvUNkLrFmddQZFMPQLzwWTsc+EYjAnDP0LOsBAdeN1+LPZe18stZ3L6AA1xpffad
8sssyaSZvaoIorbni0tRUrCEHpEOwuO7q7lAP48fuMUwQojfpveST5W/EgVJGZDgFRDJrOFQSiae
nrVY3GP9QvMEBYG6XxGaqpezTkNq6cJcMZfHy7bKrU2/nXjHB8IBNeiICa2WHY6z9x9QspfVlEja
ETPUNbxsTzGV0lfbhB3SUkAUtUNWj/kK8omzZDBziMA0CA7rY6GEBAJ9MzpaCSKRT+7MXdMW46wk
KZNN9+QUOtjjy5pJfmKm2/hoPKn4yfW6LJq3rQwX0yiN8FqOCSr0G5ccCf7M+me/U+lngmLS+LCj
VpaPvQNH39LRytww9HMpKpe/ze6XaWkjBQkLA4Ib2Zqpw7XfbhSEYmGYEig7q/v15vM8SZzH4QrH
MvwAi2T1G7fw8UsK1FWNiEqVkhvH2FW0V5zHYBlvBRR6ZW2KvSAR+AaVexJpW9sYwtt0GDiJvr1F
d0SuTTI9XrmTFf8iKv5mLr6i80tWoMpVZvBEqH58VCZTaa1vWCOrmHq8EdlncFdZYEQCJlA9Qc2a
Nt+/k19oPj/A+wj4fzwYtIGrUw4fnCoTpfzpz8WTiTvAAZA3j9qNisU77F2aN3u+1sVzJlrPEL5u
13LHaW7YstU8fFWlq75Rsq429t52fJOyaXv3c1SILQDp/ICoVRdcXZeI/5vbX0kKI7A95CG4Ru2A
+35uwYxa7hKMKZwjN8FaUYDkd+cP4COIxfTe1D+bC3FBYEVGBTaoajaw+UkbB/HFO18MiNQDbeYh
EYokMyoHTrNcALqsNjovSFaAKnezoRjgu9yEZMbnKQZFrZpnASEREHqts3gbehLWRuCZP6jyfbkO
jAIOiiWZ4gJQlw7/5HeIa/QL+nukgNKXqwvzxKGFnj3PO6w+1tfgKXLPc7HAXl+GoSOa7asifA5N
TH2+2HgGiB3DUQLIxIOjsWOC1bi2ghKRnOA9F6nYZkNKzgXuret8SQT4kwxaRxpkUexNf/Q/iL3L
Tg5WGOAdQsRQy49kdsl/KNeAl6Rx8zJRN47d7TXa/ke7O9TCYlpABnlwJW82kf/WCs6Ni6/+ICGq
JkL6WRqR4wA8nUicdAV3JEV3QW5IfrSlGbo6VANlkrdVECgtsz1g7MixO2vMm04thZcYZKXNwhrJ
WWhSIhOn+t8fP7C6rHV7qH2R9V7QA1PLLcH7bXWlzH5BBd+pn2n7ErPVVBAusbRw3qo/SazC9y7z
Ie+WB42VWtDMQAg2Y3tpGDCZetjma7SbsrceGqpZwrn/i9ytZQLp3PJ/mGq9eJvLGhe5bMUPxgoN
2LlqRKxkIj1Gz5x2e1RjoKR2zmmKGO5U6SY+F70JnX4M1U6gRJWbCqiqtZwgIlQHK0jYXPqBDITz
Cwt7xLhD5XwK7uUd7uL3cYL+VLedE1mIXs7ZAINgLqR6HKDlhahWTb7OW4HVW1Wey+KxE/YiTKtd
b7WqS+p7LDyeR2rshfDe7lLQrYtCTdhKF13lblMgkb+ykwvhXtTEeQwTIA6MALKmDdM39N0EMVZT
4FS8PYhaG3b8ZDYTB9Tp9wiRsvaWu6gyoCyyTXD8NRFBOXafeRtFQrmf7H2ZKhDnjJOVeL+TK4cB
lVJbhwEK6OrUxYnbgtVrmc7nOV2yf1MDebigQCgy2GZN6ApWkVQqr0pFYsjJsy3XWO7Nh/Dy0bv6
TIQId5nnsNQ4nGBbp8UZvIHcCX+nakAI6BqC63MkD1y1hlMVZFrnmWJp+PpbblolJLUfelxx74Gn
TiXVd91H9LAjQFCsFtQ1ugzmcnc8uxfr/VWAkFEHybPOEKpw1r07y2hmhvXN4E1dKDpZtQzCSjvr
bAAZ0CZ03gKGg7zz1Xg4mJzeU79/5nAaBbJyoCQLTtcGgWKPdUC0mdHpFFlXvs0KMtaS22Oa0f83
lAASIph++tUdAd3zTwy6y7twOnI+JAmPxMGjQO8Botc27Gz8aITUN1HI4G9A66132eZKwv3n7A0R
Y3qZiZLLy+b4VyJc4cbp+D2aWUS5rlKe+V0kk/9ltqphRjwELnUCUxnmTX1xvEiZ3a5ijyAEcJlS
BSDHh1tkM6SotXytc5LnGqA+jB+DeLuw4AB/macaHwKY9Zus079/CEZng68m6qXxgUxpwGfcwYly
X+zRtEEBvOyrKW8H+dTeazn7SLwJ/dU6je1LiyyqMIVJFI6cBukDwDK7ZD48PZmv568uG7A98p4e
UZmwJFHRD4/r+Kv5VDOIAZBB0tNNOfzRj1GI7SKQ1ns/6jEvQPwQRfx8Dk14AOLksVK4q5qklmoV
cKw4yKph3f7riHv+A61F4ZgNN8q66ln2vRK0BPB9Nd3wjHPXgS+NPQOQ0/pQz0mjwQZ6A+ZfAHrq
2mpTnecRU2THeEOzhf36+taP3cjUtrPiy4/ieA5cQgtvoBEkPdXijd6nQ9qgP1Ov/NjwBJ9/MMHr
nJ0IZm6Ri6/0M+m4oQjbmIkKUxETxFRkHx3MOJCmy0isGdnrMjLpGF24f4xnusulPiOD+ZNAbEXA
Oq9HYC2R/uEb7G8t/Rf/iYEhQ4p8FCNEV1sVWAXWFkPgOK+LUbXJJ5MlylGj4XGMMCGoiVLs05m7
mxMLJpB21ZbKF4+M/lEdRvm0MG3lB697udfGWdfX8q/mwEryonyNORYqBKbcADRe5vOpTpxw3QOL
5hHL+oBjKDNbQwtts0izd3QN/RuYnkbGT56rNsKy/Dy4rlf6OTNUMdmLNV/qQ5fWp2srQtlFvoRO
RsVAOk+k8XzKHhddBnRb/LUY85eQ93AmpIZzhlnIMHXpAcO+NNccNoiyU4OSGkMu409mfurPRjns
uMAfOde2nbFkCawQN6rXxjmLE8BGI90wv/5dyP+rQc2YLb9+spQVy4NKc1NvSVMqywbbeG+b8j2+
TpDL9nj2CTPB69+RN5+9kVcO2EDHRoj03l86Dc/o5M5stEC0Ihc5/DPRiwG+6AQ+egjAgIgN7tGj
TD6xijJjrj/3KM3YV+Nou0YQd8VFdbWbt20MkKGrF+SeVwr1O4PhuWsxdQixE1yoElES/Fzd8CzP
jbK9nqeQjQpn7sdAcGouu5ENSewo+t339ps2NptKg52cRBSU1VX8ivmB/8OaYfEHwDj2CSYBY2F7
+FtxgaPn6L0lwIzNv++F/vElo4fFncfY7s44SGxiypHAmzK1XVHwrSlf1+hp+ZUFORIKdUQ488OF
MuurYZ6GY4NXx0Mu6NJARcIrPBAakV9LOIsyjT/7muCZaExcFA3AnB4bG/FX24/KpFODCdk3bX4f
59UWbBPyRc/6sl688YleiXyQu26N8CtLM+oRJs1e4ku3wV7ykH+GXUeodIWM3Mm6Q4VLnBClUWKl
5FYQjMzmGHRr29Rs2wYmprixl9uX47tue1dDXIjuzGJe1jClr3I/hdq+3kW2Fr+FFv8lH4DOLrQY
MSn7nEdRNDImZ9oTqWtZawxjvzsGCfXKpeO24hwu8rC2Y4Ds+XuesPxrNUISqxUiMNLyHw4sIYoz
PEXgMuI7tCuqgaM5rzWiXrWYtuo7auCx1ZG45bAI9n5TAl8zWe2rVLt3ZgGCadRWVX7BQnSAe9J1
oxW3Fu8obWJLiYIJDh1szTNz9HKvjbBHDDe0+RpU94j+NRO1Bzr7d05f8OcqU/mvkmFJNW8UKPJd
XIUdZR4/YrGaHnFaJTI4XZ903hTi1zersNXP7woGFyhGBc2VO9DA6nrkyKhi7RMxPEvdTb5JXVxp
htFqwOkKBHge8Jf6pw35w6xrcLjQ0oN1Nl8vWwrR1TFWdQcxwsypXbwCXOZKcVyMxfy9suvWRuOd
sym2W8SfInHfRa8HV5J+4c9wdIUfWUJEv9PvaAL2fi+ZQe9eYPNl9tN63IwGA9UvY833KVGnxKz5
aGLbakeMhaEKy0XXlQludjUmcKwew9sojgypGjmHfuHMQhGHTxhOMmnyKYxWrSBS8p0knDi7YDFi
UFJLbp65R84+JWgfXfyeQAX3ZQoGEpjIQ6Z/MQadyZ0RM4ah37XsP9bFhX3o9/6TP5GYRFG2MEbp
ifrP48F8ajqtOytOw7Tib2QyxcAWFr2tgK1Ak68YWXO7xhVE5asYqOH1dhD7IYbOy2Da7MhGTCuh
mDdQX6hs7bFkc3xbv9RTP1qa2q+EDJsDp3QmZufBVesEYec1YR2AwZDRyDEn15qNBapOYRc64NZB
U7p7oPEG1apeH8x2ojU52CMysxNPDprxb14OpTc5X26+CozJXTvVahH3W12/yvhJoYJdx0n6Tmy6
bkg26OvqjZjZMNhmIlw0vwGMymYnbB+UinA5uu79RuNX0ghYvEjjL7vkniOA6oVgrCLqTTF99HQA
teY6ppv2qvNa9ZU7EDtpnI9TPbZkMMjkTGw/3I6E8cynCnawI3FyP4Jrzr+fxzgHR8RppXKVvcVH
uvGe99NwjTNaOovDqs12ubg41QbxojyqvDwj/bBVgC1sLNyakaDxDxDEphqAiYnM3uHwFjnPtl/9
gFIy9wX9tiAmSvluikZRyVttx5GgdUMV+0yPCgSt5iR3+K+bkdxtjr6bnIzT7u36TvenQBarFxeX
e7kswuwmKWNQplh8BnNeWu1T2ecH5C1bPfS4KhBdwLcN9SyaIY/dfpPPT0gjgRnyjzbMqLmYY7xk
nTov4MmnanAm27MTy774h3wiYraLGVC0nVFjrF1rBFwdEfBumwPrcNUm8MaJpKpS+DUEjSRX0Rg1
XWlCfLNqHn1tEpNT1fSkHPjP6gbqtBvMm/Vkq8RDFFZq3N59JYEvDRpHOQX+JXHUeN/fgUuiXk2H
WYRI8mQZRISQX1s1vQixyiqYX5SVU7KpG2X+nohhy1j09AfgoDKcm9NQel08Sla5roHHKPV5dwMH
zwk4lqJCGQaFfj4gXOryt1A/80981gSkfKCp7kIcLfJidgB67/SP63+6GLzD0PbSyCGQXCUBx70C
G3V2zmPTj/kacucF4aYMj070MH/0NpMABT4wlp55QnZfk5gLNTCXjUZ6XeyY03NDYGI5yrfbqMgl
iuFJaN4svr08kwMGUknMAIxbUEwPOwErrNukc1hUkJpycTmCiXkR7YCIfsyMOYYrH8hRCRqgBGBQ
I0F0h93jyBkCaYq7v/vkyX4Nf5Ge1cQaxreLMphNZ19XhUFJ4EEr6doe7pkW6iFcII9zE/iZUuOs
KiGUS+8mCwChdR34VQwDcuMTVRhDn7wIuzz2XhW6dyfKKdGDjIdyhviwTaorMA2f5aeh7Yx9yZR3
AImkmZzt+HLR3kuGM1duqunwbLpzzq2GNVu/6qOpupTdFXPRm4qdjztKzYS8U/1ilEiWAm1ycnPi
L5rhm4XeP1GOaCZEBmSp2+SNLuvnv0R9zjHm7u237UJ1maZoSJJHacUuWrtCZpmXpr4CdUlY4U4A
V71A83UNDnAjMAfFGUCMDms+u8JdU1kdkL7YN0mMAJ7u7stFsZ+iPb0fo6IFX6CSK8AtWTx4SUc2
YJMRaL2/s3/46WK9jDapPulLgTEVjUlKnfnLQKmd/dj99nQtZomIVoo/+KXFWfQOUOQHwkobYl4B
1b9eMHoJUYFTvbsOlVxM5YOMIv0xX6tG8t3VtZJEFKYJoC5hlihdZ5G0R2fYOQM+JKoObhNEg9IE
ak6vtcjTeWx2O9ebGJ9UAYVmeHFG5okJslv1mA2pCQXcFaYeP8T3qV2qZGyrj6oTdf1vuJAqIXIW
yObF4T8C3z7LwCzSKOH1wlFrbpmemdJ+F9mpohCfYxb7GouHpGQKJZReV9kDjiRBdGwHIm6nidBt
3cEIHV/xD+EF6EGfugbLVg3r/4Ye0XOF57k5YTFDIELfD/s5i8bhS1FvgnYk0SBEa3tpFtlRvrXE
sSil6uFAsmPPsd/GPfTZd2XgvEPDcf3KWmAwppxmbD8Dz66abaeD/DvCcxqe9QKaYeBbDa5Zo+pE
mgq4KuRz9G0meyS/g4or8fg92YWII+9ufWoatG5BR1hMj1GSMikYV+UZ4q8TkeflW0BqBp1LY0dY
qFNJRUZra2YtL0wNssRSZo5tnH6w5ASWm7p8c9QWk+e5aFNpyoSTLP59R9PzhrQCrtInkl0vRe3t
iVzf6hnUKZvRX4EZvrXGUq9bQqEwTvGI+BkInRPGhgiUX+e1eu0+N1ITThNlLC5jnQW44bXURTKf
J2z7Dxte/EkhKlF6ePvyUmxKT/A7gpRwA506WkuDdjCJpazqPBFYckV2ACZQO7JtYrip4P238lxu
ObP20WF7t6zTK/RUYITAorqerkDNzNp/Ob4HmnfpJ0Vck4k6SgkIRwxpktB8jw+iY9Tcbo0TPReb
6aHGyUErKJDeP3H9sv38CGG7qmpmSI5ZY75tvWLfDISHdSJHn2+AjnwNkv3nQ9uagX1Vh6CY1+wU
HvSX9Z0PcGx1nEq18BmAfLXzJ7GojySgjnvx3hyZ/+DsMhvwmeAomwN1AK63xV+nBVeriX2jiI44
VnfbtsZh+Jva4UZan8cQAG96Tl4Vz9v2kypH62AzksLNd7+dzb5d4/DIU+3CnRx+FcFL/svBzwtS
TjgWQcXTnPIF0SBP1LIdDO2S312+OO6EmrTnNPTEFKGNxGNhSFcmqh4dMIFMFVqTnM87zyzpnm3F
ZLHC1bjXBcMUx4XWNa948B3ZkSiqmalc/JiS1d4ndvRFcy6hq60dg2Ehi2prAvbueFoE+qVkT5BN
AIJ0SXbzznCfOWGaCilbPbL/u/d2onxkHsyE4DyZFEx3iL7xGspmtPcFo8eEYmaiypguFE3up65S
jUH6DbFfmUzPo8+5B6YdytqGLc4ahoBOB2prqcsQl8eY3BmyZzxI6BMU5dCNrSs5bRnoUa1IZkBe
uyfuHh/N2RdB9OXVHvzB9T65iWvmO6/gAVHnLDjrY+bpwgRKQ1/ceDW7wD1ngXiPRhgl/Wmf0jJJ
3ks9Sk3JrCFnU9wWbjcpbnw0dxgJYYzfiQZreyq3tWvFfhGKa2DmBgBqyvKbG4l+1LBBLhapRyvg
ntytjsZ1qHBxs/eW5b45Ng+IRhivpNdtSJ+H6ZlU4omPFozJFnQh9l5h6NPHRyrQ+T9HL+3057nQ
gBkK+6phs1xac76ohTEs229mDkVCwOycOBddPe50gpbc5gqZ9rTFqUeDh0/GyJFm9yPamNKk2cRr
prSbCgFnbXoacODu466XLEsYhllhfWo2S4hIqrE02/asPclxPEfxWpk6ZPGu0iuMGoj0pZeOV2Im
6Bb0bkSuLleazPx2W1oANYmC+nR5t6XWrdHMkmHFxSzMwpHAhuVlx8YkoSkj34R5g2HSSg/ifuPz
74Zza8ABMgKdHYjh2/NJaOb2ix8Musk2QRA8cpmObozt/T2yxUpGN/kLXAAql+6AoUuxYPYsIvr2
BkEH5jCz590v+vDgfx5gwBgsvbHjmiUsLUZnESMFLEF4+7SximM0NfJa6uAgUJwnno/QGrnYaGEo
bHoHSsx6jwrtD7eYfSv9L4DQ8we9bPD2iwavaMepErM5+Gk6u1hoenwOvYBYcu701x9Mik6brFi/
iFzJZnKb9TSREJaAvakdB97ckelod3FxAfHvEKvwC3q1GR0Xfhic6GSgjn2/tSAz0Oy4u4IBzruK
gcSRFgwKOuGI/KbaZQ26VKnLJOWO8+oLv7CCujcwZKEvby8PoH58Rv8s67SnnhocV8eMltzUtXhe
vcRl6R9ObdV15dHKHTBQjhPxT3LMbdIEwoKeeMagLYkj7UUaDIJllxyrmyuNgrUhMzC514RNC49y
WkyyjlTVH2FcYQq+lAd8pVKneAPOYGFP6cpZ9JNjsM+VRTvyxM/W4bBBQOiN+hW17/3vgxj2Kix9
G3LcxC8SdAahb3TBHY+D2OchlsGm9M911ucwhjAW+DNr9vDC5+L/VOjSnsDwvys7VeLQeYTuK3qh
tlhzzxVWihTiQ7/eOJpKYR5XJI1PQCvxOcGozkLTgLzgZ5I9rdBE3KSrDe8G69omXdPgUdqMe9Rw
08kcvOKiS01gzt0xPmSOxVHtNqO8R1kH1JTP+nmHVyAqZLQwj/VNDRKOiJbF0fDTPPSthSVWBiQ2
DcCy84PhZAeltZV2a7ZO7ks9sfE3j+j4Uyuh3+2dExxW6JE+KWguQqXwl9oOfsTKLlZSQJSdjg8x
a+VjAhS4X8HEg7I8krwhaNdoDlsHIk2er8TPU3NIIlWYrw314+eVchF8fy4kNh+3dNeIu4NLri7J
3cgdB8nov9WYNwNc+lgxRiWTrZvogCPCuke5ab1lQLbOtBjv9eu4r3S3uYxN3XqdaSdNEFbIk1/l
oRk0L0crlQKRA43G2TQevNNXiUW5VwPfKocivAewHNM33faRDfWGWPbHZf7d3/SmZW7h7AFuEe4Z
7MuYVz6pkfMSmxCneoKjM0xU/CmPkd20n+0t0IcpfO/MhtdRWzRSM0BzoUjsQ5EGVVUVfO7J/MVh
ddB6eJz5PKXpHTX4QqutFCBjOFMpxW2qf/y/0mNZfs3laKTNbz+W1rT1ng7V9QcWsafjvFA+dT5W
c+vpzV535AOZa1YlH442gfwKjaJdvRlPOoosfQ7JTbbEgYBnUfGKns7H3QgCzjnCanu31YkVittc
P5fehdlS02J+6ldlId61aijRvruZubVp/XwjJhDQb7CKRJ6Umc2cmYfYMB+smZyVyPZf4IxAAt/S
vqULi9sjJXjFyfm89+/L3q6msTqhIlJfkp4hfGmuo+kEm6Xc/ih7l7fapf2xNi/6xAAcZM9jKxa1
zzJXyC5RaUE7UkKGxqBp5h3pj234hINqZQVBNRFvIsVeueUyvop6JLkvZxZRmvVtgbrvGJEbliw8
uAWMQ94E8ID0MvkNBev0krzY9A08dWiudeAlD0KxtTS3/czfz3iYc8X9oX3IqAJQ4v+Jh8i8N0Tp
4begD41AQeN0YRhUUSzcOwSJUImU7MGUMyUtOXbsOr1O0CFAue0yzUJvdrEeW5/hfaCdSptgpf9X
0c4Okyb9cIFrwkX3TV1fj97JgDFEP0xgblObpI058L+zQyaBB41et1wvrCKn93AfdAAulQxBe6aC
AxGfH18h5n1BE9ohE52WU9LXsU2XpWjsfN93ibDL5q2MRXM7GQrByA3sNVdG9KJ9v5YIXQoIGDmK
TBZuAaBCqJRo65tieIpTWstl5LURzWIu7bTG4K9zADvlicKZA37z/fp4SnzBofgL8XKLATcphiM3
PMmgfh0+shHy6vROOs9K1QoAVtEmhbrL4x7V6bMLPQmeoBGvYThvK1TEyMUHB7ALOpOFR8aYriS6
9Q/Bi2FgiWRUepH7xO6anSM2WNZ7mkmR8EY8RMTUDEZEmArWerOGw9ChbxN/pWna4ZHg/Ru0PJWm
IRwUhoiI8xctcDF68BQ3q72OZAlCmUSPTjw8pp50Wh3FqjFhMhDgrzOWiXiVqYBZNMEJj20z0Hoo
xpkfevZjNu91oe6WyJljs7HqUOuM4nvNPUiPpedCD8Rs2gYNNHnkNT8eO8mzfNHWSCJoD6RAmCv4
ho4QZFzVqCHKdCIoNgJiAL3DnkOfWcGXNWBzAGlWCxRewYBWGd1VjoPp1fI17OXwXIM2LcMn/8wu
zeoEJBSdtEqwKbGf5JwtGJOCA7cptMPE2JJmU+VKvt3aF3gkG51DtVWp+/xu8qiRLNTFYwaNYegS
jjV9VRUq8wBI0lJ8B5yk62gr6CldWhwIrYnlwrjoNnHzby5KLreDos0gJHTQwt4vGMaJwQw591/C
zXwlIT28/kdjfnXmxFqvmbn8Wg278l53UvxNHYZh3lG2nGsPHUOz4bVGrF4ltDK3y/86ApGnXwVt
h/Po6sMceyLin6rpHb856JI/9UMn8s3piZYnlQwoFjrepaizYSBL3WabgZl6uzsCde49bEOS6zd7
GuOLSkARKzlnjpQUdTsXhl40c/L8aduiHHs6u3D55bnnuncQU7pzEA1JKYL65fyMXBzVRYhvX7px
V2t1AL1GROHCBeL3/MdYozlOQo+b/RKoB7O0MIT6ddXgqMctpke2v9FBcDuKBZuON9twkLE51T4W
EMGjY/JZmqCJPwFN7PPAHQmw9qvO8nQJ9VccsScMZacGVZxAR2zI0kEIrUZ9nOD+a6AjEkeXWSvz
eXlPUw+7Zejm/wBZddxdOuQF2L6VUhDkrD8Q7yaz54gxCAQhzGDmGjtdc06CYOWYfqoZknOYipsq
JZysuOVV8n152zOp/YXyczrYZC0vJHRNHs1g+VegHGiSlDNbSFJuCjJoCMbP4qJJVIxe8mCTmIKu
ljYz0CVfCCD+drgAon5LomrAgJBzpGOzgoDobOHnMD9AgH4LZNQBv+BxVMzjrSoAZ+FlktON5t9D
oTX8lDFyxvLpbmSdcYQiLERjQCBFB+Hi5k3eOwKGi9Gk12RfoCnjjoVbmTnXDVbIsfGRVw2xIHxe
UzcaBoB+/N40W7saneoHt6jxDMqceLADFeM/0Uv/K+5tNHFFqID7t0y9c2SBYWWVUNQj0UCxW31k
0XVUNMxemx+n7C7xTs4xK4zsyGxcywbsjJKw6jY6Flylq2Qh2cMN9gKj/4mJhBguCHTAZK5BCG1f
SDxYBDYuflksS2yOXQKq4uIUhUY5zLUPxLQjC4mehJo+qpusDw9Qn/Evj0NSqPjyX3IWn822fQJt
1AONFECSqCRDVOq5Q+j2DA+ygcQIa2TjABacDtDKsm2DcySvV5F+IlKDipsmFasVN6XkwW7MzUqZ
gkAl57WflhEHswLxeQdwWCHea+UPGD2FkV5/wuzC0u5BuFL3Z6x8pAc+NDf7aW3ae9BfJPfPYH/H
EC3LMpqkp5wCA0wrMfIDFBruxtuvwnyCXoNfIYOLgTRJqXlUwMdN5rYd013ZS1YN7pjOwxCATNNZ
DyDptkr4TKPPyZpA6vh6TCYJ5RQdM0gygsdYvKB9Vbvp15w05v6J210k2IfX0whXuDqG+RvCY+PX
rDNHkvzxI/g95otc/x5x3RSotfEWmu+/DkEDBFm4xTDd2QLq1qRo3KStoYhDOQvHfGHnO7e7RKe2
DWsn1MTqfzohRrswXwrjHZ5VR984uKRI1kDT+jHBo6KnZCqY6fqr2p2j5nLokPZ2DZZkJDKhv/1t
SKKJcN2ID0ArGSn+6C/2ApEnpbDR7taF1+qu/kRh7nctF8wxk4sX5dKQl1B9xGhAufBjOc4p5HgC
9//ESIxwEy/dZQGO8vxZXDUO9bkq8R01+0RSLbJCHpKtQTxjcbeelCgnYPR/tgXF9NguDIX2208g
i4ml59IfqrlVaZMQqStlwaTZz2+4BeNK+TgCYYMkmjBjpQ8lGFvWo4MHE2IMXWKf3dtzNZ1GqOL4
pR9m9ft1N87pU1K7z+wHeXub3ZnbSQvUh693DFU0MfZpDBGcBk5Kj/gy8BQJ0slhSgvvHQVPAkIu
0xUEr9g/THWB3ZMoUR3k8ZyNovGwc42l6NZkD2QydDH6F2XN1VaJ6woTZH+ZW79AzuV8rll651/p
HXuPtzZEAofp25itB6cBLJm5w45CWZkzbjTWQnaZGgW5g+DxZKLfvu32d2Pj+oC2l9LspybTpf8L
ZFp/GdVrT1zujIMqgaeRBXajUqj+1tNgA6kdhRNUOVQ8569RrwH6BpeBNdxABib3RIP2e/htFphC
7CbmZrO0MdkCz+IyWMQDEeDTedHs+W7mIFSPcCG1wlMjysUN9R1EpFF3p6cw4F31ohUdlEh7lvGj
Dhq/1DQ6I+dhHruNeJfvPMHn3ikNqMJJWyPmAfx/lccj2tEFpm8vq0KRfxaSMUCwIWdjp44nFvFR
nCcyph2eMlDFf5eBd30X4kamciqLJXEprVx44jxQbVQglT0vIeKV+x62RfPy/pmonQy9VChw7FBo
Fjl6hlNeLDQEYne/UA2ewFtd5APAc1jG5susGNpZp8hDLNxHFaPEM2yyRf9TN+Qgs4/ccgwNxL3x
dEH8vGfT3r4qbRkdEqDYluK7tLzKNzKoG979+1ZUCPs1e7sbaP+1FI5JLDug95dP58JfXSpBlMVy
/jJAUZcQOoQAnwhagtSizEI373QbVnf2JLV8e+E1316tWwXTYvzW3UzLaMvZCuYB2UsO3fpCXRaZ
/1TraaXgOwg7FV2TwjL8QI4+51ba76Da4kZFOwl7IglckJBUdw6DieoVWQUFvBqfP7xwwm2vyrCY
Swma0FCZtTfa+P1uuQEDs1MeesE6M73pYQVz/kqOIE5OAmCp++KVwmdQRlSVhR4D1vyqDSJfNmDa
TF00kYUD7b1mg7WU9s8l84hdLyGZnC3gx89enrzthpmvSw6Ywp5oMs3h0EvPjkLanDy16n3CH+be
BivQ0+SjSbQk+N9dMnq+WNGaBosSeLarsnwAQ7bPUMbtux4dL+HT4C1j8dDmPj87nn1fy48TMUFj
WSYI/9gFP5NFFR9+y31QQEO/PhZYZaG2wDQsnpPsG15/I8OxN7U9KgQLcP8U62XkkhWWpQyIpdGy
eXbr1Zp8X273+yFCK35VIdMONHK1qeAnIK3zQp82p28Ko7UplSIo2YFtV9ll166tVsXztWNBt9x6
5erpAdRTsYn6z3/dQHQg11O6feReuon1Q7hjoscKoh+sSFRhzI5AkpcimeTk/Vh7ZVuBQ7KSVhLN
Pm09e1n36jqz/ezYz9YvrixDUUK/KRCGdlSjCZnRiLZRAe2p1pKu69jzJX5QlFrLC+n7CEx62itD
xPpP+IwH/ytrReypj80srcm/Kwl6cLl5bkXO2s9uejIjqwPboCiRhijwaB7DuiSpwotDk5ArNIZu
qii9ABSNV2XEbenYyfuCLS3Qvis09Z20fRsEI4nJo7XvIQ9kHw5Q0mUEx7D085/OjIUAiq9Z3lhJ
mNkXXkPPZlavZ2CbORZ1nlDAett4YUJE+LbuN9MuT4hpOPm3xZ/4oD/T6/k/hn3KR4Y7/SPHyRne
06fTYmmp48KrZkaAVFQmOu5W+CA808kiygYIGAuyg4eVZDw/Y2+4oisbLi0rXXMiSJQerIfZQ1tu
fqF9v0JfXIuRQQriW6ZqAcWMmuHNLXotU2dTo2AOmpexw+Q65nWl0CpQ1V3ZlAVeIZPjToNih9As
wetgCx/04HlxY8H8ya0SPejh7PtSGpI6mJSKAvBA6jfKxGDgctpZ9/vpjF9rnU9+4cSiJcCWHVAZ
TYpFioKZsXMGLFi6rTpZ1EvQu2FBa5+KB9wssZeAhHtZ8z2m+By6r/RXFmngMvQKtp2F0LKcghth
8ga+B/+J9HeM2hyuswAus1IeLGaTLj9j0rxM29HELrdTNBzoOBpp2WH5yqGNEko3gjgvjR/4ZCkl
2Q7VTzbtoOt3RW6wR6yTNmy9DtENu/pA2Y+MsmxDf/IGy3O73dCZDOY32y9glBziUqpVLpRY4r8J
8tm13qtREL1/Yn4qgdhWSY1CTT2ava1gVjsPliVztKjEh7gVyhnAdSbkr+zUcVfnam4FdUnQdXql
rEwbdjJcxZLZLnbgC/PGX67FX/rcP7TmsSPLRlWLP4R6maewsTvUbWMIYr3WQolF1pPMrgoUyunF
OU7UnQVwhtPXtBHTXtA0tGa3MekMKebxG8yn+GxHXmbrhlji0jCZJPo/F9KwdwT3iy6HLlj4YjHo
YahSr/nX0zsGksiHofDamBF/+5pkdh7ipGkWVsZaW8/vHQy315KK0T/nB5zrCQkWTIX7BvUCuq6H
ESIDoMmqmRWYanA7uITlTdHF2Jzyb6kHpIle/Roj2K9PKQsmlnbSqhF2d3jyXVIBYoqwsvoILHua
bJ4ptQizR6pzcV163Jm8C8A6PAAC6hBSCq8Kc/lJlB+8oqdlkYFMsX0oV1Ej5VSt6CbrriW7q8QF
dBBg0EofJXNoVQneoCCn+Pgbm2KQsjEgQ05ChhMme3+H3/onZ19gJifnJFrDH2oF/LiyMymKyk28
tAUCUzBp72+XGLIpxxq6bNyRCjfTTbVA9gnvp4s0e7yl8eRP+uRu8jG+Pn947NMznMfFZl8knR+6
wBIMaYxEzX0vmlH1bBA4EUU/J1/ciLkKsazPhRZ5fTATMh3zyZ4/YLCbJ/dGpa4V9DlUfT2rHS2r
0gADjp/ON/Umk0gKIs5nbmnEw9NN0rYvrROWuh/ZyDgfB93W1S4Lz72yQKqAM+imcgyWiupsGuLA
yO1Le5d6oeiX8YA0a/nzK4nBqUyH1lDu6sdZcqkxWbXywiKSP/+WK+YTyKj5npJBBUyMj+tfFYnZ
RGwh0GwJQZfOcmgQ2b1b9CIX+qT7n+J9507s9bdmydTR/ECNK4F5Cum83DYd3tO1LRQfCpq3ZDx+
0Fu729D+fLGufJXyxP2M5NaOn4/pTtKsOwgzEr/CHIRlfnJkvIbgliOlshifoRUsJzMLzfttqlk6
8NNef+3INB47BwlZKCvHFMsil28j4P9DCLElDIQW2xjpj1FagCPN56eTCUXNUJUbreWdFVCOg1ox
jFndVukPxOup9rcQLLULyoYV/H3qholP3RS4mUZzPQrgQxpqBP+nVPoc0XaQ7ysRzP1RH/RrAQep
rSjAiqbqolKzKKWkys0V43sMRXm7kIwcwFzh/ZVQw6dposcc63yDZKVEcsTbTPNeMatVr/vfguWu
/K++Epp5W45gYydbOWYAg/0IZpcYWyv/nyaqizMV9cNvLKszlvqaF5+dESp5JexIvMDKrxNwkUa7
6OM0CT4Y+FYIMmZGGpbsj3I2vwZw4P/GpzK8FKo2E30lYxwBqsktJ/Mz92NmEW45Zp0DmXKKEUpW
t9+YTwrnFTULjTA9i/dc7Ftp6NAkeMMO4zKiU9QDBjIKJJ/OoezHuKuoKDstFuIy3wYrHH8sFDNM
Z+Qrq01WigHitonANRwiZN92JxtMIM7TZ5sGuF/gkZjoJLDrxZ+2EnquzPHivCIQcMa0NuHoqOjW
MNHlG60zfF22vGU+NBE05pMSsq31lCcBaXDhOX3g8DWvPjTW21Q3S1+Uanp2N1D1bCHahAv+O7w+
u2+HvCTNOu1h7qDyl3H7o2Lz/0fqZZCJkzWzPcp5GpYkQ5kHTX/xTIvaTPAEKqxjmaEMkf9N1pqL
Aw6ERtaVJSMohfZheA3z+AOpgAUng8T0cT4OFnSIF538VTb4UhuJVVkWJM32anKfEJJ+lDcCS3uw
eZi/JEvX1FiAd+qIa/qWDIoOwHroU7wDdyd2LvSIv6I6VtOC8e4cvGHFEVQOFwBvI1filMJPLxwF
uaj3qKRWmu8rJJPKjdPjhBt98WuMV0MmtcxKvQA7/K8RYO8gS1Pp1xmbRJQOmIOzNL24CTgft+5N
pOsfmbTeJxa7wSGqoZ4bM/BALAXogKijoYRt4TGHOU32YVfZmxfMDh/xLlzzyqHxZifGFSZAa3Oe
eoBxvq3olDNowsnd+0YNvtPrksXscKIKX6cOkXDlS0UTCLICAe7jCF3dNJ0UkMaU4oHpg5W0DirB
gKx9IaU7BfkYqcGCR43Ji73EF4+ZFivNdEqRP2RZVjZI+9JQjEnkBMDqXqiP4bNJbQyeyPFKvZY3
barmtGqgpWbRYu46TK6RxHdCgNLx+UPGeM9CUGagYCAvFEyq8IaIycPVDJYtQUTrXFMwasmH8NCe
802v/X4NnT0Hkqvh7NpEJESlF4Ebrw5BhuGvPaFIdDNKJPhseJHPbaPcRe+z/lw5zqxkZLBjqElK
lHvOftTRsAOavFsdZjBlpvfIv1mNtc066YFdZ7G/RoHOuDkf6WD4OzRdpJh3MPmwk44S6zJ3ErXn
A/LW6HouhwrlGx5zW7tdjmDI6PBbm7N7/gOv8YbFeijSUnIw2ZTTKhp0GDn2vqDWpPBprN/OP3us
ZT56SY/Ejz4m9Jp6NQBqD8JS5VsEwwagRt3RfihUrlqhsOZPtP1ZqDmZrMeDQVOLTRE/+E5N/li3
WLUyG0jLxpGSBelK/7mX58TW2po8I9zu6RnCEcTVb7MwbArnzqdim7XOfioGokAnvxRxxegOhU1O
bpfdHfuy7kzjh2g4iC34skNJa1uz0ba41xvhf70vumYOX2smC4gglHskkPSxc4DWRBYRFsagcIMx
f23+ySF7DTfn3A9NeUnl5GVJZecPuoTGoTt4ZCuT+QXgWVc9poCvdXp0f5ZUW48udNtSc7nFOw+g
JMrdvlcFJ6QWMbS8nLg6s7MMZkgDSx3T07s1mYDQ6VWQD1nQ2z7iPKhkJtGegkrVIn8Ghh8ypZFq
bEO0lOr5+mGnsoWOGGm3a9GC/FTIp/hu9kaBqXCH/6ExXQ8mpLyMkNoHG7FBLC220TCzuhbbvKdm
83/Y5rXo67CF0SboIRqpjpcFY0NiJCyU9b2qcGRONj5QkOKy4GdU0NOvHs7QlM/E+gv2f+03ABgW
GTAvPY4KJU3E+WNpEvTTffPdWnWRiLzCEb5e5ryHrJzq7fHbzVp/3T9b+6WcxbfLGS2ByRNVddSc
PqJzfRv6joqBzcwJ7AAusvfX8qh6+c3ArzGtDHap8JgBBVvnEFRrKLO/FQA6kZCzVVDxHQMrcevR
zOJRkTq/FGM9QJdHmLGYNmTlSkcgFPKjQ/oH2UEF+ijpQvhGSgb86sXWhobksWPRwGzOQPwTv9Y3
sfK+E6YhV7o5YrHDlaO6Qn2FoEGZ0nbPKzxbib9uGiFGcsMZQMLdqrZcQQJEf0vDRwSLo4V3zjF6
YuXO1sYb947d/Avuy6szG6hqU14CAOGsV3ry3r5JGEQnI5iKV+1XdOo5hAKKyXpkXld461V3aVtG
KcDl7/QKUI7HElzJkVdV/TtEfvcpVae+EknbsjEoz57LeeN3w1QkkTln9m+F+oLBw/BaH7Xz5Uac
2BaAuwZzS3L2ATzvl3L/0AFz2DNENMBDa6WRR79eHxHHmzwnht+j5WWloU2bLCG8tEZFrrgnT8gn
h6cDpighdS60rIiBSMd65akFiqA2aM+Tvak3lEmuSQixVQhTNxKaQKXI9b5aZxb2bESxPR1RzR96
9aB80+53NjlgogdoLb7rDYViI0oFkf0vAzU9FPHn4/pJ7l3XkJI4c8R7qmWvZWwFY1XRSmhcRPSl
XXKAgNazrSEfVqcgcOat3Nr+J+rANCcYOrDM+gxuzPWsa5tvHNHI/XOezAGuCbiuFUEBzDxiQFDA
acgKK6Yb85bGz3CuS/peU7W3Ud/S2ZJNPF2G+b1mcVypX2RiZuGUwlv33zepAGcJvdZqI/13kWnt
ogXuVPdjUJsn0igI4gLK9mDnckkogQOnQANQrYxYIE99UXsn7nE9kSZYrgj6hCYokDw2c8ywpO9B
0BJe9z9oi2wnfDo6WmKvPRq4mJCEHfDNGlSM55rg12phpLicwYgXTPtZLuu91fr5A3RaNqGmOsc+
/XVgQUNGM6bXDrp88bMr+u8sICXxVBb1+Hjs1nFJR7u3Lu1F16hjX1cR7YFC4bQpQi/nKPGbGOsT
IS2Qqyi9cAAxMQnu+Fw2SzHkjgIyl+xwMe8xxC7O//J6fNvShOTUU//K1lKZHKPHKlPQTPaBkQy6
5Nes4TMp567NB+SldZmxSsTI9yvP4gONuO5S75N9sCExUt5leLR1yxAJQ3fkCYgy7YvAYM23r5eR
89D6VsbDdc6DZpzJZnsg8WbAPtkFvDpqObuLBF5Q9hy40Vr1zy2KUZa+orNs6bm0kEGWxdmsQ4VU
q5vf19tjPykpAsqDzD0IO6Bi01psgQXVxRA7QSziAjbQOBQ1jTfuvztkGHg1QJ7u4q7MPqtCoh5A
4CSfx6vhuLTxmyz7Uw7c0gDXUbBliooLaMvhV3mWBox2xc4u1XBhQz/EFCSJUd8Dcl5SvVExnvAf
BsOHUruvyUNrNsVEdVQv0pek4D6UqVqxHWDot/uJrlq9bZ7NK6x1f2BMYIAK7hnQoeBUfQovrDRS
DvaAp0VGfmAF4HcXgXyPgyLrIHK1KJP2/BleYvY/Upz/m0R/ms9SjUrfPS5BqysxiF8wxi4YQ9vO
MBA3eaU46PZyxcg5n0NjjNJRTnRZLDmY2l/oHLnjP1oT7ANZHTakQH8AKQgeBOtmhxkaCQVVU8zM
OX4dgfQS/Sxc8cpXoPOXSzsiLM2O+qrppeK93Qc6VW94WkNRrrl4vCy6taAgoVgpdRf5i+qDulsh
yKKtneDpLXjy/MwWw3xY2XF7mwt0j+IeuRbaNaLVR4B3+gPTddSPgUrYK8O1/fZ5UN8A8m+YcFKW
tJf71lITwuQXcVh4zTFalPxjWYNyJO9jJrGJ48L6wY0aEi3IsUn5xmqrfT6QJfrGAUkLL/SpBleA
NHfp1E/7fK63V1wtqTK+Al+mwS6AWzSnIXAu5Y8rI91JYVoyGexbQvU0aDWn344CVjFl48jdkQLp
jL1Hk7HHMsLP+kxLWhO0743mBoEsDR+L+oreGG542U2jyZrTlnNVAZ7+ECm+ODhqpgTGjZi+UR7h
DpPAtIjLXV7LSSuITnlGGo6lpNGRTc0rKbf6BjUI+cP11cwUP0nkpr/yDo1h7HfTz1fs+4lwRKdW
Z8pFJymZvRjkORyWVjBncb73UtVOjWW7lo2Pd9No2LuSNtVIH9Tzb5SLg43abojt/dP5iI5cQ3Pf
acMI9KCnTGKedr0x82vWhtYi4nLah8GFhwHphPJL8RrS+eAZKsjs0lvLZfno+2LVWVzm8tpUcVVs
/+lwBuAxXqvxUbluyEVr3dRLoCbIEvuvEFjnPTI3hzxlq78Rjw888X6apgFTn5qxJie2p5HbVeUJ
NRb8pLFDXf6XeQh1i7i/qr5QjXypqTffYDkUr/P7YWRjhM1QUaXqyh5POFAeQovcFyYMenLpnirP
yqRhUJuSfRDNE4XDJcGQPu56vMoKcDKJU3WZQeFf3Z0f5HiHNg5v1F0BzD/J/ZASuU/xx63yJ5vd
W6zCt+bLKQIhrMqn08ppTFBkVhJiejVWLCMGbT3bCEHdHzWm999lCnLMjWBuNneFsK7D41AYeC3n
LW1E2O89C1vmrm/zJyoHeztmdBRH/3m5vEbY28tGedxZvQiGZW0dT0cP01zRcAJDBRbo/MV3Mdtd
RJ6XN/LtGEoYRo8U5ONjMXO9WDkuPo1MZIeCy/7/Oil1m3YPZDbDYXgkHOq+KXd7rya3EqNNwsE3
koviBqdTTlcj3XsG7L6L6must1c4PoTY0u/62MTT6wg1aggoQ9autHCY3pihaszSP3jojKhSHJPC
3MOaBNfbihVeDGdCrVnmM8nbyufPqgdXsATM8buoPaKZ4BMEoBCXMuz6067iJINdvZ2cs0wiFzq2
huCP0neu2oT1A/NcmhJxsxmchQvGpWX6VLDhUM9Yd4mfufktPC5kX1On3cNznK0McF9YjnWTGm0S
HJpG5lFxvb1WcDJZJ9parQUFG8IsuT+8MXaLctVI21ZNOQ5SnmYn/tGiPBPqIncY/P4vswm92A9M
9HZiNUxBwbmHji4guARn3iuWDiRsPixShdbOS+J/vV7CrEDdKcuJaDlyevU0oQ8r3CKLe+fk8MK6
dDWMNt02t/OuO3IUSY62S3bC9N1U9AILHJgbFdsLXOubx3fYTJKmbttgNHKGUxl24+cX82grEnIK
F4BKB9Z7va+x/QCBFfo1XLHBDzIRm4ROVtI+fs6mcD/8XLG6ITC7KTwGN88VqDfcv87E64jMXPKp
OZLH++keJ+65NnmtPRP5X3a42wwTYiF5aPjcA5VzQa2VXEuwNjSh4IXGX4jB1pprToWMRFn9R8iY
FJPyVxjR1Qnry6J5dXr1Yoj2J3reGDZZko8002mr+8frtBNuDl9gSmWPM46sGQ9mwt24fGTi6zit
cfWo5k1orpqRwQuRLMkW1TW3d6YM2xonJUSSZyETax2t1NhvQ7862Ypq/3pz5A+rtj8h6SFuWris
KYCB26B52VYo6wzGD7lUbPDzSCwiyafUCt/abnagq5PGEKOiFiHa2wuLOZgYo0SgHPkix16ftmd0
N3datZwdZlk5nMoeDF0H5bOutzeOsewpX4vhaC+mRtXHk3pVjJhUprYmtu+8XKNwIzsol5ikaYK+
hE578yzJsKnJBb8+/jQjGMRY9H9EKZG/wS2BctehANxlxc0/qH68pcIwpScaYEfNgbzgWc3rNzEH
AGMkr13Sx7w5FTp89V7/0dbVgTpieFmXbmUDRGD1a2NaUHUTvkzQ57A21L8MkQNt+XZJXbYfa3wR
tSAy1ehMwKN8OAfx+lMjfD4frngWaBocuKsKe74Ne7PWpjKbLH/aQX8nUX4iH4qhLDO+9gd22/bk
595iaZMvkbvtPeFw0Tk8heI9Cy6NCEbc75gpozyeYyXaxARaBN10K0eimZxZN3zjjPJZ54GtH5L7
Owx8WFmQ8qF55PqSrxIwKyFFcOOMuaO2eN19eMeR1WeszyMlUGOWNuq4Dky1Baxng35P8lx+e8a3
IT1ABbhKidiQhVFH9VZ3sEZe/pKtzZTqCVdh/0XiMGwoX7tOkzLrSHsJoNNqkbjTsIs5ZiYb6Lu2
hwsmID9nVIasEyypyeN5Bkj/9jiBdKJiiUyOtwWY5N3WEOU+wUlWrq2qIVsglSD2KsHTKnhcmVRb
sPzOnHgNurMiGLUzk/4qHKOqJ8d+XpcPIeFmQzZ17WKpxpliUCMym0AnAaHLens6VoxWg1jRX4xT
v+Bl07gNFMjS45XwxEI3YfSND1dVvS7voktwsqiNy0WMLrcBt3VGNHHZM5xpf4pGfz8iXRXRwZVs
tN+dEfx9gxW5qyzp5/SYgD+ailVpa3XOng9ZKjkkle19h7SJtU6FlyQcr6wxgV1AxRF6CGx2toXq
V0FBrFa53J8IAskGfGxAHzQ7e6c3DN+KGFMDcGsGlyGdqQ39RIlFvN9J+s27GJrEvyjtiAIqJUCs
gBYOLq+IBgKSRmIFA/PUDvLWCK+odUwQ27AOYseFuTzVRev35/JdIaWef7O6+/NWWBMN2aOe4aYb
yepPwThBEqa5ONJkK03I+NRUnj5TK9CgkzuD4NmpFSaFqHz2Imvv0PjVHq2HQN9qyGwl6hlkth/a
KS+xNw1z0x/VK95C6sRTIg0NfWfSxoICFQ6iNibArmg1oBmVUaKn+/iy3t5TNck4D0YLDrwVJUa2
Q+IPrtMhmx461B2kKs+nUetllT3ZU51oCIjRX1tnWnwP5iuvFzB6I1n8rBaahtLdePEXKKGKosvn
9hTRC8VKuouZFdxjFbRz4gqGd8wGYwubAVEpuU/qWm0id2rb3cDCeedSYYJ5wHxdTRH6ZJnYGDnM
zVrpo6kDXlb+56VSYgyX4f8buYJ0NDwgqf/5LtKrSRuXVauMC+eJDQXNdHd20aPqmczHLPznK3D3
DKhvJoVSqzDnztlKfhNWmKEtGgZHjrf77EP0nRNi7LQ2G4wSvmr1M6tAZh4765lAC7pVvI7YFSfn
58nmk5fGrwRgM+odeFqV8bOoenoRp/J3/gdlkML6hqig4cyFwnlpnEDy5UHmXsQuokxGEqlotgpf
wMJgYsMLEhvGKdMl9FFbvZu27eaTNtBQZ0oDhiN8EPeeHMPLbNCUl0c353zgwU19nxNmtAqCYxUM
vS3BZxMkLuIW5oS3Mtf18qQNnxPBF+MCnnkZzT5a1Rdo1ryXvTt4alHhGO1dIM5+0sury2GOGJIF
/0HQQ0KYM1rR1Hjkg6bmwiAgASoLiBbxDQeJOreN4esinzOOjlz9AwnIjw/+yeoTMT+wDO+5px2S
XVMaRTHBNNuNIED2c8J4MXDuTtL4UrxRK77Kb1yExMGHkzeFfrKvAQznxQc9g+KRpLBqzFD66GvJ
P+LFaRDIwpmYMEfzWhpTMRYs9ykwperu04ZtakQJGceAnjo8I9w+fVJ9if5LhczxddV+Q8vRVdc9
+l0WjqfQJqrSbcMkY0vRKcn6XZt0IJgyLuxTRN+wt4uRey35RxXJBCe/RTEXcfB3ziyhfJqpN1Wh
c2T42d2ymJ3ALizcqzt64bdoAPBDt1IUs41RX5/RSoUdl9g2bShy38IV+B77NDvW7QXmCPVBxAqn
22ocqXx+nxbsbtWJfmIfIL7mGOSyN72vJ+9JHUXjRccnhdgYIEoMKVnqqa1g8g97ANJ4nBmA5sKW
4UwbUl++WnwfEME3HG3p8ASoNyBMAUElbnNBz9lmXroTyY0lHfH0LxxMfWjQjzdhoR1EuRGYUkg2
by3BKos9irDTEdP9RuBQL2OTqSe4QBAFjmIsSNdLxlgFjCnjeWHdtX+A/82pY0sFjotjZR9+yVZ+
XhFVxHz0dbuj9DAE5dfgJlEqCohINY8ZzmxmfK5A0Rj/HeEAus/NpjmMrhpLr0knypFRj1mDUtPA
ARK9tvHyda1JLkoEwawLKpXwjkwNFJ6S84sDk/KTPcHWadovg5hEQ2c8Bc/HCzJATHoFGvO7fxrc
2FGyWHjOzOTXFAsrL9kwrMo3u26S0AgSczrtik+KfJFYXSiosjsYocspnGWDmRl2gk/Vbg3z4Uvq
SunZBB5N0CG9ji7Mfkbgkg9Qi+IrKZtStIxecNtoKLqPDgpn2DwwVIu6Y6BoQOOM2RtCgh1FCzXo
DCb+YoVNRAdDdfEcyaAthA4oqqb/iKa0OjkHqBpfMrZxaQR8ooTmgkjV9Lk12AT2PnUkxyCiRxyT
MTVTo3kO1phSHwS8C+AZ/fSiJArVf9PlwOyDD0KrQypvg9VKKuis931KfAclysjFuO3EUhko3GUQ
duO/dMMZVEEZ7esR13gNbUhtE/BXg/XiEFB6r7tej2REE8fyS08WknXgm84xTSVJ6K4uL/h4RIpW
5CNQNp4TBaI6bn/i15lyok6RLT3QzYjqIPDKG7Vp6D/j5CSO209ASeOQRUrIXkcnBbsu4Bjmro83
fwaCCIUfGiL1ZlV/YG/zJStq4ScZ/oR8aPyRVbfllwtkxU/CMjP/Yu6nkMlji/Wp2qHF61kO9+TJ
OSapArOzXYiP1A1r8a7vAUhnayIQXz2kWHa/J/TDBQerWzeBPYGG6E71ak4Mq4N6ohRP393ezvVW
9kB8eN9Zydym5nx5+7TELvdNU/euFomNGLMixOD5qkDCxqL8AJD5MwRofgy8ZK9DADhym2zx8Pit
Si2Uf1ytH6C4ACPMsBWxH1yfEwRgRyOG3DTcFYsl4PUAV4pI2pWG2MSRcYbxd4fdxwKctlo+iPIz
AM1F9XNZwQM6N4R58DOQU2PqV3cYNhoOWgQARUcBubFjqmXShFqSsmxGcBl4XLZQVAeCqsjxZymB
pQt92SbxUcnDDGh4mnmZjHoAf6Q8GHzqpzJriU0D7F/5IMhVaS3yU6ltloOjU9I16xoHHlhwCIx4
vNxjzrQc31jdUN8nSsqJ6k/RQQb6l2fLRkBy/MiLtrTCM/Xd1TwMYgAxv/oEXC/OPxQs4EULv7ZW
Iz4pbTfVAdKPVEuOq1LAZWUcvMZPAG0XYEY9/dbYDymzBoxGcBdG7t6OzxyJZBwuD9Jcf7IazC6R
InbzNGY5xQP8kbOHW+QmG1yl/p8mQbtxascP1xsHwrlixhz2Q0vjj77ztDXzVGOEbfrhskb0meYl
IQKfYaa+6WxgvLEzPnb0syiTXP1nrZZJE3yctMFpnodIE0uPwDyrvbEgfUGo3KB8xtquLewcAuq6
7+ieaEpwzBZRdgMXN5DeEw09YO92ZVQaO19w3glyMoH5ero678Vztt2fUmH4lsTn5SdLuRe0zmH7
kr6YVE4nm/UtCa23EMrDKAYfB0SpW4flumHX8bVWa/BT46zx0IxJQej4xBdjmkCu15CIY7dqy4vl
WHcyWpqIHsR2M2t2qsMkY5tInN78gZeUZBUot7qbM/bldq7TXx8+UBVlBeMYIm7BwMdM23x04Iih
IZdUzlguRZzcmERHPZFSoMJN6KMdRr9ge5RyhbRSZHW+j/01p+ITd2fQsghWJ/QMkpoqXJkZz01N
9VsnnWr1PjRjCmcoRKvIir51rKhHMlaYg3TRLvb391LPDQkomS6G0iRVvDkAivCe5c9L+jjZJgTN
SQMV/X+MeLb3u05Mldx10NqPj/oRozcxPrpx+kbk+69CpUKlI5FjsSh2OdiKJdCWSGcr90sTsLbF
bHtMEs4QVvB2JF7W2gI8DhL9A6R7ayGqzufXZCYSXmjkoyZPW+ArrfH92cgMf+t4FurLvmT8b5cw
iu69UB9ki5zp70AqPCmqgHR0+BviLdJlg1XjvfHye3XafLMoaT7IDPcti0AIg6nQQTxmdrbEw8dM
JId0MQwJkQNEVbKz5G78DOR8MGHduTNvdoRo0o+bBOfqiXSTeQMKUTNaVKfOJHS728FPBvAxYHBI
J0h56a8GSUEkiY5UehXE9p7tqjQ/1h10HrWm905bvQdtLHPerJ7tKybvFk0XoAmHfG6UoPhqh1YV
II00mJRvK0YOP8MKYiOQDCvoomA4RrY5DdA4NpejKgwLKOW78J5Hc3lfdFgMyE4vWJbOOILEIFZA
d8XENjmL8fj2T3bO5CzXI8/AF1CVO4ao/wZr4vXxGFa8aNMvBLtlmbDQxsoa1uJEYpAGcytEFkxh
fK0FNnZIjFp1m7N9zGlJ+luNyoB66Wtc8iqPRM0D/4Rd23Qc+C3sapNzGZsn6fhX2HDFkWUfDzvu
1MYeR6yehR2qnSvVFKfrHDakWzHx0AGXiWRKxtvPqWtcPcvp9Nd9B4m6U9NBJl9D+C+LcuDYNmCC
Ko+zjtW0V4/8nq/9n94JUKtO6Muj6TqL+p/nJJIuJNq2kkBaTKBglosB9iWCcMAaEg720TXP/VJf
J/dMJedASxR92+Oa/xnFjOuCIvpOm47fawJQVF2qgMyau2tNGXZovDb+w+nvJoMgTCGRcKI/H8Pc
+XF8q3uIjnvQzS66myLycXHcNbGhLhdL9bWUkPengzwUp2A/4YJgSNwJrHsrG6lm0OIkybdX+HaB
jI34XTfrPRuz5pwry3irIXCSYul3SjFzxN1BuGG1mOEYMhnPEOUknArCOSO9bk2HEindRX31EIC5
Nsa2oM3067ffHJiudmhr1X1IA3yd8XmRLS6o1bxm80+1uSihH6E0w4y/B+p0dxyyA+R3Z6z0FXza
lUjY9lhi43b+O+ZqSOSKZ2j5LUFy3h1JYdM3xr/FMp3UBPzx7cMhZ6KnZ18OEH5EQM22xhXMPfun
66JdroRnzv7cyePAcRTgtd9ITeN7JmTPYzXsNaYNRGbaAxSytu4+NdHilRZ98jpMY12qXO5c+OZu
ldgy0PjCY+h0Hq99YTrqyCYLUyDYXTsNRaUt0OO/qgdK4xWdwoxq9bQqNWYMjLusHvHMpmR8J0lN
11pV2MSjaAS8/WXNmHE9rtC0aIsbQG264edBfdaIPxsq9TQqCGXgpSLdORAT/vF/mFyJunOzSL6J
xVKjurT0ZwQrQhDlqxWc9ZSBIGSn9oHTnf5VNJ4wC9Z4VLH5F8tJgs6fCssN7QuQLhhClkX3usZp
eHbX3pt9kh/mQt6+ruPrsACCmq2aR8rbFYSXtR/wn7RkNuLE26xVWREmuPyhWUlG2bQp0e57Pyw8
fNeiYf0e5wZ0nL4mA5jVN1A9fEh08EMz1pCM1MF/CzInppqbjkhNSbPM74q7nMBpAZl2hXyLhkXg
/U4VdQCPT/j1Kq96Bpy84zBIfyAmHhGBAkUwJwFQgocnpnMxCntpb362Xia0UiDKrTcm9gDsvLYR
RZ3JUDnN4FcFn3uU4wBvqCGhRiR3I9LA6yVAD8cmTv2TVWSo2/MD0VlvrTTNR1m6HyD+ap7okwDm
5MmbN6cLLRqcd1drFH+ZoY7IJx6akX7B5xt4s4/KEDMk4jh5FpYw/y245cmmgMs85Zr53ShFCcQ9
3blWThmwWpjH09Q03i2S8i5WkVrsdfHqjpR0JnK6W4+eZGDlXmPZOiqKwhzMf/5BukRWv1sL/K5D
bU3JfLGCYpFDbke2xUw2v4zJeW/Z+CqXeDyNch+TrCmWf5qq9z+AR1pK0jEAWCZ3gEWpsGR8xdzO
7T60qh4JCdAHNJ2sZF11SRCvZ4hJh44l0ixoXPJ5utFJ8/RxMZWfRSEA11D48z2+/8wgFdHdIiBQ
Qz6KIf5UNrzdNAtw+y2Hn/I2po6Sfr3eGXeiA8k/30YEjpWFoUIOjMln+ujabNnADYFdIN2pECC3
NFtcSfO40pnLn/mnGWfucgkMBpiS78BNfVFwDPWb5UMzrODZT7eHHSeH7WjZ45msWqoO9UgVPL3L
/k+mI0pWiJq/SvJRqrdjPZn1StUYBa4h9k6qLkOSMcDxpiy2hSaD1aRVhp3npUeyyNOWoRsLvmIL
Qv89OSnVO7jvIAx4bX0drQG9H9M2QEzfzHd24N91jnoHaHIZ7PhLYs54tY4Ohze1ILYQ6StwsKIh
m7pR5YxW1e3VRN/ckvqzq29aJTcp7B3/q/O4CcVGmAdUX99Ow3CmXhaWsAkd+OFUaF1vl5XzeocO
vgFKT53O7GfxhNzM5/6QmwEJskxfNtb+gCCP7kwH2in3IjELb5uzjrAX/63LHYBf7M/ejvrzXldQ
xcLgmvfxtF5Whmrjr/tvsYzQClh7V7IfjPyLivhRjVRo2ajHobzQBPN5RgGG35iHXSHOCepKCjq2
Cp9eNN2nb++RQ5C0Vnj6Y/ZQBDQXDe6XJjlMaq5KzbQW9HTOeKnfu3hS4qDecZEEDZMwYmH/u9rx
FBnRA99RhMehGH8KFOMGykLwkwMPEzvNhJRyvu4nV9sFHw8Xxm6A/X3aIMU2PqvLb+ZPFv1ciaiZ
3sv09PDA/jdOJNWyZxV4GlAfpX6gL/p72HHeX//+hVV7tMDKDqQIS7LAWMtYKd0nzskAxKgSqWQ6
KW7oJqkV1wQ9RrU0/BKA7pGcfSl0hlitVTADZ90SPTzYpWw7Yj7CCapiHow1FjedsnM9lDEA7k2W
/72vCkBJkObieIV3ReRsiOmVLCTuj2r4JZlvqPFzMqPkgOWQxwselOYmLFmwfxOVIi1EuLSigBbZ
3Y3lT+0M/qTSuSRF5eVZgu0oNTF3JZFT9Xf7eGzlfjTWwOoiLV7PxJ8Cpi0p3G41jKGWManpEN7k
AYaK6XTACCgPMVYRXCJyLjUiESRkFLp3350GzQpxkSDp0FnbRTNCiZTtdMZQkyOFHMCWlKvWOS/3
mfrNEf2KRWq5vxibQ2ZwQdpkGt4fo4Z6Iz2/91xSGLy/YKfytMFzsYgNeXqN0mLRDWrCJyUEUkoN
1HO/Gx9oTK/7cMGpF6Pj+xmCGsobOLoZsiycvg88rF4vaMhTnX7OesI5wUxVpwwtKVxS3CrUEQZU
tSBZEwwxX5HKz8sppiEbBaskXUrzAMw/jAkCibc2zmYtMXCZKTShd05HylIF3wDwI2Hu/XfslNBM
NUyeFdY9On4fgvG2uFCOq5J0DXbKzF+WT9PJfSizGhgr72JMUhEUOt7nx+he4ZQb+c/Gaby3vPfm
bY55TcCMKjpF3RfNZ/BXhXJ5wQoBDAXOWvjokfzldouC5Sr21wBWedfITuMA/o/v9cJMI2smQSt/
wC+vTO+chFaJ196w5GA3aHK8hFbAfcuODhkX8ZHRm3QDiE0Hst4nqEyAq6KZvGHvR5F9HNtjMwOH
qbNrBNdDVagJFjL9lV4TBQl4B8wZfGGRk504TdoIwRQweJ3vI+axH5sMEMs7tyDGT45i72FZ4wBI
A7n17Ag61w4ul9tvAGcGSsEv0I8XGL+ebPpdTvSNfSk9AtsVprihG3J3FLFNRHjBaAXyZ2WEsNNl
mpu8A2DYYl8VcUnUnKweoJoIZ7fp54PxHPoujvz77aW+PHcJXLek6dmEm9fO+iBbOI9LbjYu5bOb
6vAl+880tLYgAhs9/jk5FrQRpiJPBmNIjHiTEefrlzTg9L77l31+mzrPwKzchww1DG03y4ktXR/M
l8sH6f/OJioWAhMqDo1bRxSprqVb1HpmZAzd2DgarRYXz15pcg+X1/ALNXY8qKHA9GSy8cL0Kbol
GRSU4KTs9223hQavBlTxv6i7G2/xlWWSoTfSnr57Ti4eFRDBlAQ6tAsRNj8pMbPMi4Au/hIvmfmx
ZcVWaunkM4GWbNqeMEP8Jznp356w2vP1O5CC1cZ5T6ah8betCbDO5INxR1NCR5yjbYDNSuvPNjJv
GbXqO/vr074Y6Fx7iAwCCiCe4YORt9R2TCIb1zAByte2Oi1vahI1Pa+aQp8y5f2LU7UrdnSGVGUY
tB4NDoR/OSLZ/uIWZN2AAaFw6dLVKCWnID/gKyY0EeA/4ZoaTLVXARJdhWDsiE3xefHhXw+1SJO+
ePKHxurrNJYlIiBdJk8bBb5rWAhN3O/BozFlcPlJUXJhJlZqw5zRzsmhhaJ6wQyTvFJWuCJgWpzZ
LLCDYBNgLIeWxnk8zIBCB1K25vykMSQiFznh++tz1MLAdDBYhTbPeNg5FETdkPDr/iZGXwYMfaa1
v6GIX0HGhh+I5SUc5GW3iVCIDtSgFPbJ7wgMVK2WtKCVfppLBoXm47L0sCo8izDQxmu9J+Z6JQH3
wozLQgEswrODmDHBWKr3yPgA9GH6ODEQi0ljuP7vLeIgX4ftTA+xCTva2nGDJBr5NiQJJIZNlAnL
7GoDgMqZc/ohLQ2GsLWZUUZKUBz18DbHdJSfvtFQv0IqI2Jzq/VHEp1ut841o8v2ZmXxUnea/hLC
VOgwPmwlsqU4OwOseZU+h/Ztt6ovwn7Y/jEJt6pyk4Q+R3IYYqZqWvJHwWogUj5GEgPwBwJ23qvV
nR6EZ7W2xeUuNiVUSnfadX4H69XRu11GLbVAm/V+BhlZJcxct5t9YgWn7e/M01pWb+hNGmzjNriq
WF4BLrdRU4hsWzLTBMLu4hnKa6tv3V3vuQ2NhSqI+H6DqPtSISAw47Xlc5q9eRKmHtUcFLfNPLDQ
RKTBlPwNLjPfzP6zwQGub5O70fr6APaqLCTcNN+9bIOq85iLBtw2RZOfqRoHbRm3XxYml/7ZqaMr
GJ2deqKmkPLOcDTE+aEBYmAxuCNZB3S/bs3F99W4eFNKr8RtQIVpEPbKeocgzGP+UDIaohJcd/yc
xVCkyGsmQM8UewTNiVl/yccHZuGCqTtQIBf2/NjQkSr6JhOBoSrHzUUt9PusnpU9rvEep0KBQvfL
KV9mZIWgFo2p85qjbFQT60Mz6rN6Sj6b0FT/jDGwNtGs+4Veju6n71PausW2hJtvQA7fhT2Nk/3W
uo3ytNpzy7GFe+E0T6i9EBXzOJbokBopXk2Y9EfDaOx5xepR/8jVRUTlIPzm1KSM5WjriNTuujx5
1Ju0ayeKGvtjv4baSIV6nfMAD/VqbyesYoEr4fA7/a80WfMgvhKUv2zPcUa6RY0OjJQo7PR2Ire5
fCN5KjDVL7OxKsJeMKyI0bGBz/8VOxtPCajpVxYIF0PE0znkBJlb6ySpDmL4W2ySyr+PQj/3XBrC
Apqqa5Yown7Las1AmZqruYO6MIvyxAH3a/PMMltDixsPEOAbJBeCHw17OKcZXyho7RakmCEr4F/g
Wu7U+wBqeUX40hDu/TLjWiu3z6NW82ngITYXdeu+Q1nwxo4PsX1zkjILNFhfMfCfUqv94S7JwgZt
RzmkjoJGtsvfXCDkYF/7uOarMhRjjP5sSQbrrf0FuZDzmhU6KHZq2d4wlkbhKRWQz4Ou7uu+27Zz
Pjn/PYkOLDMQtmdjd6aZdCDRGxyyT8o/yIvv1vj5Qp9R0Upr01EQRyAyuqtb/5vlk+PNnxruFaWi
Ft6GLeBVH+CIW3QILJ5TenpiXnxtXc0IUAdiWcVl8GNQxddNnZzcIa9mIMljMj1166T/rcX54lTQ
Zj8UQGcYusqqohVfXog5Cc0bsCZzjWxZymESsB2s5GPv6RNOROd92sVNsbf6FgxFBUF/DQ7MjTaV
NVRucpteVHsn/y0DEghjiJSnbA4m6SfJMoPQjTp7HL0YtotK92S9ocj94BxQTZdHTU4FQKWrkFTU
Kqq0/FotyC7OAJgOix8Ur3qTgojI0yng+gxtq7h+ZhEevpQQHPT90R8DnAQGrrxXub4eKJbfb5uk
kGtzEVQzBhDZLCLfDC83Ni5MCBiQu2VTk9m591KmE6cNjVFLseAIL5gGftE0AA/E9H/SDO2WA0jD
R9UNLp/5YfGpNusFeVxldPoFYeoakvJYHK/9Cf1jpzYGOU+NjisnXrXjBFUmGoZEdSmRn288cFpW
qNdXPywkQyHQBTZKq2ETPISVcU6mKvZonzAe38SLdMpTeYPF45mflcyFaxmzgDp6ZZrNwZ4heiAc
F6+qHNrNE4a8cQ8f6eUnVNOTeHGqnCjgcSf9RXmePDwxwZKCUWQovTzPSku0Zy5lYGdimSzPZlhf
58fgJN8kZCkh+Mg4RLjOMACw+IP222RCE44Wr+231Jxaw421N+Mc1VsLEffvdL3TKzw9Vj4jN9Va
gCb/W3wSB5TvQv4kZpavZlcF0rtQ0QYmHL4CKlLdRmmBBGrq/z/rt6Gt78Cx8j+R2rytnOW8eJ8e
Rq0kr6HtN3CvNDnKOq6TBt+6u68dAgjdqdDc6gcfqOW+wvNPt909UhjCVwKrGU0oe+ljIo0oTLTC
Ez+R4B7yzaQiRnY4At98SBPHK8yIjKj3SZt7bSCnoIjyVJ3a2b6nBYVql4dxGeeISgaeCxG3AH8i
ex/nSddFMh5VQ5Q99EOVr18JfrVh0C4LwFvQTpUyVQEmPAR8k0d+yJL8RQgKWNpMtDml2LD9yKLP
BWG51n5OeKDQvvMc+/F0bZ3uigtJbm6Ae3mSU4ygiQPszWUvj9+1sI2N08Wgh6jJtDSFv4O+os+q
Ffu+bnkNrvfuHhNiDl0jqx8qG+yuiUuJl4konCHxlnPk+6lLPnRwgIXT7sLSZXf1283XKR1qjkM/
Af8bbcPG3jbRbo8z2KHvJTo8Ytk22FupGDCyNSsJd+3swbDRpeQaegRfDGwfhiDlpKgnVt6dfIBA
TZlCpb85MCgoMGiTJQjhIIwiol5v4TTNZcHi2kXYsUy6Yh9r2e5IsYdbKkumFPcchyLq9btfXZfA
dj+rx21DfnSmPBHq/a02w/hQEcFx/fR6k1zD5X8pyTeXpz1ilE0Zo59+mNnl3BDuH8grsEcKdM2G
2hkokLoPLoigrLYIPfWsyb3StWBq3MIJuv8vTDJ6xXjZ6KTA0+VzBphCczUyscq4V1BpwOCz+z8y
PIkwcxTAWLEHli+jalc7bBXdHv2jalGM8BB/ABXOboJAyisNxfOletIo4IYVXsMv372sxJ14R36z
/EIQ1gjt1/uCnn+Rx+rVBnXkX2HKKOZZvQIZ1vxUOtx+T4aJ4a2UMZFsv+cON5332+7cjdttEX7E
gsZWJgtiei0BCCqEmU6qryyxM0ZYIvHOS4IGfrq2F/dqA9ilbFqaFfKs5K3bp35PNWOiq6izndXl
BDNIvk+iqfrq6Yj7drG1k53HyMtcjQ5zJDP8FZD+JsCagnGgDr+nBX4bqIN5h+EgF4vNgidCXCB9
Izfotu7rNtyU5VzZ/Gx5P/JS0BonHUN42I8EOx82HgaXWhc2ZXhc4kHHQyJ8fKnVeTceeTdN2WQi
vTTwmNJetgQ1Q6izAMphevwu6E5+xj6GAzVp1zGP7bcRcXeuSwNZTIP4jgYLRjbZBeV4q/xjLeC0
/ZNiEkVvzRkUiNifOOMgJWZtZBJjyGLQBKdqfzb3ni7T4meVtvQDadnN/CM0xk8BkJReFLwBfC9N
sC7I/tITc1wlIRwnzfNzt9k8KHzSgiemcyDZ2NKC5nFZEXcWvBi2OLUnQlvkOzNk5zXKDJxW9kaP
7xjS+V++z+B4whrZtnQudkhZCS+aCprydKrE8ClTR9AvXs4wtnLYDJST55wY8LLTggRxp6JdRNd/
1wiTxGlpWNsbYEZEGE9t6CAl8ndcUKYgu/VkDXQIpYxed5QVUM+2RFIGTCVjVCYV1ZbDpN6ZrvQp
xgvxuVfiBIUr47WF9jAaFY59mVLqXd0+MJATSfAdZjiDi+dw4ji5YsSo8sSi59aTmJYNOAvS7rKK
znwj7I6g29PRny73zudzJbAIR70OC5B6mhuUgIGz15NcMC9TWYV+pdzZtyWgkgu4NjkhKn5Oa5+1
nwoaOZaRYzdeftC6kE2Jj6kNSTZH2V3iKvX3ZkEOGcWULw769TrIbWYODf17zv2eDfx9KsNC/ZZC
Y1sy8wqGMiBP2aCIBQgD+eEeMU37p7v4GmRx89ii7uueFbXi+NKEX14W7kPAUn7k9WqAGzn4fIcc
z2NiNENT0hSo+0WMDA3G2q9CRFpQQgFnYNJiuAuuDgDrj66IRctbaIcz0mLnBE3RIahTK3TlL3LD
FVY6ZCSmdQrH96QTYh3TmDzwmBYdPrseyVLKj7ayEci0yvKNxqILiKtBbssN6FLRrgSydJsWlyjK
AY0xVXyKJ5Td5lQJ4a85p5qlFCZlCFFCpAcTPbJB852LZZm39WUQFWvg31H6/UnBZtZ67hzu25T9
YDaVg5jG+X5j1RGcdPFh2J3pXNn7goll4bMiMNltFIxfdKD8xbfifIxSXRPMokZvclmRdXc/q3QI
ydUvOQtE0hfEwbVc8XCrd8wKn0X2i3yiQowRndyR8Uvxu+Wi4zp1G09QF2kkVSGUfFsUTVOeMhVS
bha1jOtqE0L2KUyd+BB9nMO8ci69xkNYzVuZdmU/1bC853WpnnCds5k0Vr3BB6pkAigF4XXrsjLr
NIsYrSoyJJN2TW87d3Nw0UgzfoVSH4/AZPnqDcmDOaB4AB2gp+NDUZGQGi0cikIvmMesVwwTb7HB
PhkpH3fbQRqWZlvg9GEDONo4qMUiLBI/kff8m8yEP0AI3fbI8QgPP+dlOmEi/iTDk4whwpVzFkaL
pGwVkH25fG2OsS1HK5zzGeHNhcryeZ8cpw6SokChqj9zkzNgmwPvnNHNGplrktHnZnarcAhIogix
3BocU9CONAxp8njOeX709cNzNWioXj//0E7OS8jCpXTDnqWd3cv6Jg5fwdC9oMTEjQZN+kHngBVz
P+L2gtoJfTiENOE1rJ+nNa4psnyrB1pVzPlE/93G1DOC8UbYPfss+cQ0hEFTJOb9Xa+bBIuYOdH4
iMy/SsstJ6ePFgDSgOzZtMl9AB33MHohyJqKjAVtdHVsBx+dXJtqYNDvRcnUfKcDvhWOB4U0o9No
BBajgB72/XnOvpGWu2QaXcb12INBJ0pa5LlhqytUtAPWTSWp5bdq6WTBGSCSm3m3MrBAlPJgnUNK
oSIzqlXEbBj7no1tOScO5bVV7Ay33vRiBqBWPIMONqfmUgKCQCNjaP/D3OwJVC5octWOLw7kLQtA
mUbLFJz2ceYlrVs+swbX10del2D30mw3MbP0fa6xdOJ+MBwFXTinVOthOaEHVx06rk465quNGso/
OgpRe3Dd0dmWPQ/Tg7ffdr79689QX0OiIWQsNo6y8JKOa9qgq0YE/yhyvlEQYe+5Si1Qjt+fah6D
iYRyqYIPIFVVGATyIaiMKmamwNV/XpqHgqKFuajDpCh2ELK156IiXKXI3E5r1gCBO93h0R7gZnqE
ODTAVMuvsv8CjJ1cc/66Sv+Z2vfr81Z+22kk1bD99/Z/c7HwoiMwZH5rzI99+IbEX7gauZS6hoML
Vq94iCJu4Z/yiZVf5jREBANUjKsm5GJZNo/6gFveGSnK1ofa5AAeGpcpNbtuLqLwUzkginJ48eab
C2sq1lCM5rlLvPtPcfDt/5rFXPHIUn5dRp8GmbbPZ5bTTW2vtvBTUFKNY0SAQRGYeX9pu48XAIZY
Bzgbu0QvloOYvFLE/SGKbeb8mh8sptsESAMbmTGvBn4ATwut9zK6Mg6Zu060YSZlNfPvP+LoBmxV
f0qYm/nBex8C4Yf2Pnj4olFb6wI6n8lnj98FQtQkQ/Dp1tJ1OU6chPc9kFJAU84w8keVtKr9UDYd
bm1ZO6WerHtqrUmwreKn30rAkwgcijnHx/TbFFo/sUo1/aE0cT+guXgKdrZrU1a82pzteEro6eqr
X1Mx+NID47FVvlMTgq3p8QVRroEIy3KKauQZgBZ8cBvi6Lcvpu8bvK3YFluVrawijqa1GuLsaF2y
RKsQvLRiPRo/kli0WV8I3b0WheN0lz/B4LVqyWhT+sawGC5ff4q+ddUt/qoPI+m7Ygy9n+YX94/J
TYDvlpCdvAt/2wzCFSVHg+JkXGP6disL3fFUfDvOkJFZoNpjC/LGWZXsGJghJWlQXRukMwht4Y5l
Dta8Up/Lkg3JrQWLuWwrix+KpPoJ1qAH1jw71uNSrLuXUHg1E+B1UyLtwmdjW/t14pjXUt7lzRmd
bRSwLlV16rlRqu6wquctvIOGYWLMh2BuHXAsc2x2a2SxVkqBVp2Y0yylSr2bdyIl51eNXXWVOiMH
Wh0H4Hw1rakfYhO+YRKmQfVdawpSEFQaVQWF4vPjQkml3Jaj/sg93my9mzFqQ/5qlweBSuILADa7
tmZtjV2QXhpc0iQJsgNGQ8V7WYQ85KQMbW7NmbwouyvOxhH4/d2Mr0d1B5okRZOWuXdVFmcYkxDb
ACud5wDuog6I4wage+xoSu6I6b75b7cWECOnjtt+ygNaLApQO2RunDqqhkya6ubN8B9lwoJsxsDT
MKjpGykNNPnhIYcc3wckyv4Xj9GETcrGNbZQsP9xEUM3yYskHXl2Sr8TpYGp8xURkbw0CyiXABja
JT0fOZTLfjy6xjogVcTo37MTHHEA2/AsyMfBkGuYEpGwgFKzH+rlx34AcYQcuLY5Z8OhtIAcbADm
cTLUrHp7MI6YvGaCRNU2nACbO7CWN0jB14Lo1V6AEJidDkP85oFPevtdveemWcdxcIH6mTM6/DW7
uTtMPQNI7eLh97BJaMPpCm14io2/9igqgnC+qwBB2CGQgH8VKmdRtcCed/nakpzrsxXR/0DFfau3
LuyurdfO/EnZp6THxQ3GDfeNHx7WrPy5vTWNlweCmqlToWzc3nCeW+Gufp2QzLCs6VBxHGpWqZe+
vJRunz0LSWON2KQwwLSEeZfwXgIwNlcvCWma8xvB3DXswQXAOAYrmbr0KoZmtToQKeCXVhf2irTA
4sV68JkoV4+IM9IXpYkYTzQVC51i1oWnHkOHkmpa3Ni4K+T8krUIoC2A8C7Qmkr2PvonYEAzuKn6
MC25HMWldwr8Y/yJNDwMr4M355/+SfPFj+prwE46APQsvoYJLQGhR1jYZZuEhrnPHYTtXI+tYU0S
4GGxqu7iSPCCQHMWZ0p6wBmVWd1GF9s+m/GR4KapkKC887hvFRPu2zrfrfCXULyiFEkQw1Jil0CK
veseTR6MkzyKj3ivseuiVgnoNV1nas0NLTVJmu+vBBKJO4wP+zqnXJlFAKj2+GZz/u0ugpsAoJe9
Q/uxAzFTLH0/VrHmLjR/PNpG3PIia7Y3JQoz+vH9+ekqISY9ln8Edx0YYcbrB1dRIo5F1VsqHBwe
406Q9CM+zVNdJDrLQs+lZlasY/w3H8B646CIWnJYC6aNlIeU9gsG64s7B5ulESPbdRtbHx6j1TX6
TqbxHsgBbi1U+Kzc0RAS0r8qmKqfwZWtuLJdsVQ8Ak20nCYvuUswuQxjvcpoSYENLN0neaX2V634
jThz+5Vyx+AGYIGBVMwkmylfwQY5+6tyIWwdn9xKh6dAxMt73q95ZZGkIhBeEMen6+W6UlK96bti
YaSazqoGAXCC+EojNVQgWRaXDPUTa8oKh7j+9EsPmmuOPcQBH0GPni/m9ZzX3z/qOvEFfghxo+vq
1gCo5FGk3EbVR6yqbTy1VKdhyMseS6CTg4mpWw9IaqdqhAeFcDRQjdRoTMtk2KP9pz36Uayb7zQA
0r8C64oAg1Np4L7UDls4WJbPFCeMh3CrISVOuJW73HxDlBdmC6Z7XellYRKjzUH+DoT88HZUk0Db
LrHon6Ut+7G911th/2mUl5Zq+2DgQ/svKvprrjfSQfsaoQ6FTv5QE1WuvlA6Ya86M/tfIruZ22GS
1dasbH/wbYXdfuw77cPvvwqYRqNO9mgLGgtbFtvloIvjluN16xqPY8mE8U4JCtwSavRgQPQxgK7F
L2h4tpl+XMEblN6lK5Ig8R7qaZ23I+3fTT9gitItpueKozGLdJdWGj0eb8PRNegnzv/f/ATDH8eU
+MiOfnAXK+ZuXvpa1cUIZ63efDGrdk4zHx1uYoqDwbgO0ErtmtWfeJy6ttsCnfLvvXhq+LlvVYtb
piRt6vN+1uj5kjODRCNyKfLXaWHovbM98PupILa+zmGs0oXuIUAuc51dOjlfS/QyjIIP5JuQUMwG
kjGfhju+xu6vP2ygEaAcIzKagwU8sNY/9TNkjP+XvHkoYdYkX6TiCYACSxaaA7M+l5f7TxHr1sen
CW5SwMuoHRa/DHBJN+fMZNr/gzVypVWlNFwVSdb89eOqaZeQ2mw8EQWC16kK7QfNIpGRXRvKiS0x
Hb6zmA2y8Jno+SNhYg0SOztxQWKn6pheshKDqcVj1O5kPcpqXw02LwnzeUOjvLLjQ6BcVWhgeTZi
RJuzKqHJMOSoKnDHv1gsJLz5vYeh1NRPi9auXH9Bt0jxRtCBDZm1UBPLusKPRLx3eQBA1jA9qgyj
QooF4olOOOAfrJFbwIKjoIBOuZsZMPJCIAvyVEDUhWueiTDOa8kdjKTmH9y5OlJ+Wq95lRPKqvvc
MC2ldo4duG1GAVBx5Xrh4zTnoQ+4L5bwP0g1yUuRzORgtjsWTHF1nC3aHxZPN+jRx+4hmsrFX+R4
bnhOxWCg+ZxAmS/iFRqxH5LrUHHtmC8abInP7aisiO5xFZlIboVjd1c7nUNxVORdkE5eEEa7rbce
0Xa+/qABH8g4wiSCox9RK/1lkjUDE5/RA2uVvhJHkBoiwqtL1MgiKW6eyz1+LTd89Odu+thPAYVc
dX38+U6FXgFlOcrL88/rLN+B7929YDkPgX8D6R45SK2gvnZBg6kEFHkNFR8zWzXiMmBSdZ+6uF4V
wYwlUYPU0WR0TtvWwgD2yUFUqEcIdDVsONGBQ2RfhTyECZ4Zpj0XQJljPKouTsfpd6JuB86v49+E
xFV//m4pzDiAlIbNvavTAmMSRitx6dHpQ3xGsPU0Xridy4oeWmtJWTOhVY0u2o6Q2aqtiXJbSOsk
ntKYK6XjM7A5fis1vInou1u69Lzjqci3PFClg6Q9IlL+qrr9rZETr2gKgFmpedhaUSOVUQshqqqm
UBOIbBVQQoRex0YMoXKqWXzJrwnsJ/+lUrowDfZSVRHHRVp05/lVC0sXFOX7OygtnxuRWrgd8HXb
1gai74K6OS10v8agl+FJ670GZvMCAPhDrrD10xVdQvoqXDRHk8kXpvtewPkXcc+VbM2i8Cnuh8Pd
96qtWmKz7+46KRQMCA4jwxFaHgfu8QO/9ap80L3x/duAxOiuNw694f2ZVGlSdDfzddEp1B7AS5gl
T1+CbI4UVDaEH42EZMIBtCcjhGaJLiXvGhKO3+9Ql5vxK0JIJ3ldMAw1Gt1c2s0yE7VgKkgbpg8a
U3zpm9dFS+EMP49I99hBglDmpEmdADUze9sFw6NW9S6baUnRQo1M3QnYJ3FMr4L5iyri4MOMEtl3
opwLfdiPPjdIb5ZBJeFxAWyO5wvDWV7fN7Z7bITJon4vck5b01mWPoty6U89lecVfR8W2Qynu0Of
LgTbdnq39LY1ZkK4E9kErObwGnIWyehu/xAu0Cbh8lIACZqY15aezTyRNenJTo0GXQ2cCEMgKbtY
0/Gdwcg3UPgCz1d8dKCXKlxQ5mTvsYpwBQn0e8TgqyBPj5Ay04rzKz6PTK8eRPBeEFb9JFbaeFVT
EGVtomdmausKTCKSdP3Mv1gXxvcqNWhFt4SeFvGPIymjL2kojpxbNxvjNKeQUipGz2Wxkws8EQr3
3DGJCDTYAeB5NbcM/vf+mAt+oa6xb6iQMueNIUD4eJxwbeagdiXMI3H0QCu7yArmMXvbw63qFlWm
vNWyZVLFDtTKgY3Xi9ZkcXHbwTArcvloXpciXGB9ptKoe+HqY6eI4SDDqdGyXpDor4YuzsH544/x
T/XDITTd3hfRgKtqWUVrJb9d/f0SA20vLXILtJLFId0Y3fiL75OSuagH5D1ed9zQIeRO0Ir6lB0T
d8gX0LwqPp/Zp98w53TFfegLYXFoQ06CBXQp2lV29G0c5GlzPll8Xt2e8pq57ssz0uZhv5xvRcEB
mhT+5qFE6806Q7MrRne4yKabOD4aShU8NOOyMwaF/7kfhXsj8bobZShequbVRXtX2JYuTfTqxjjX
MvBNRH+rkhB2oMUdpjGYMm3m19FDbELwTrOcdxG+AhgdZcGUfOAzJxdxYBjcwfM0U2YMU4jULdTc
Q4lgydmHoqzB6Jj031GPtTADFiyDy7ro2VBwMBnwLStm0fiH4zu98FfFUHCbM305dB5AJcd6PIVm
HubzALMA795r9wE56GI32qvaCThWMgogu7Ttdw3Xz/BdD1OVWmWYwb8ueDUdN24P4Fqm+hscbHUs
zYzyD+HxvIVgAmYOlNVLKskg/RDqSuvlglPXgpkPNZ1A3mPD70P1f5axFyW2rW5YYnt8TlcCvhA0
Q3jPNJUwUHC3JGShuj0ceMgx0W9OmCwmMgp972D42C95nchDHKKGqqnaty5M9QBZKUBrp3laggQb
4JvfBmtMNjBcxy0YPRDnV/PG0LiaNqBtRsp4NtB0CV3G3i5TJlhQ33LIEyHY3SXAhv2Xe20/Nv0H
ecjOnsw12nJhcBU87rowlOz/2LiSlD1O8auFOleXMY9YOGw8KY82ZqpRfjXHPxPE27dZepLVLvaV
0swFEfDid32pVbpxYm2eK4YzmaINgrVQroDvGPT8iU0SdP3vk6hHI0lu2vQIsWh7GJSQxgvDRs94
MnK68k7fMUxMjxThM+YX2jPfu1EV6gT3V+ux00xyRz0cRyajpjrXk+hL5SZsbvBALzJ9yO/AcSM8
c8Ja4k7W+WcNombdrnXXG5j+E0N/sffBvH2jT2wXBTpMhcmRVPjPkPqOI6yvJeV0Xuwj09epxqf6
6p7+lhQP3ZEKce5pmoKuceYzlmz6s62TQb88PWEqqVJNrGlR33CZTSyJ1JbXCl91uPQJ8rRGPEu0
DkhnZVz6S0FkkkKEwODe/4P0a5DhCXF/0OI7rjwrZ2gRtsSs4RsTcTtAv26wEFydVeit423+Mw6x
0kZdZpr1EMAIiwWib5VilL5wrjmqZSHkuRGfHrgiZZfn6AH/Yc+FcxwIrbc78yNK7foplf6H86vl
loVTwI0ttQgEWsRdiJdYwu/2wF0vQ+qEz+8Y3TgdObbKvaT4sy72kzcxKcRCHZHBOlz3laCid6ld
yiQt7V7B7WWqjdcy9nYjhHcUnj2Ja6ETULaychmkmTqkUrwatU5XQLe2fLrSSl9F14HqAckUuxow
NcaZMUe1z6U2tvyug0ItoQq0OqNz/mmp7z8PNYr0gUc2WB7strniuIfchoOK88CHW+vR/NJSRdHY
ljeoCvGYKEktNPpCO2SjF4Q1OGhz96GG0c+ZtqqvoITpk1Wn0fin6AScynXO8akWUDWWmCX2fKVK
dzAht0+0QlDRoV1oB181kvvy/BEj58904eqmtDRLOAEsQmJnrQcj9k/gykwz4a/UUe7Khh+766+G
yRANuiVJdFegNm8GbShzFVrTFPrr/rsSs7NIoTfiYSFdCMUTwTj4hWkW4LvRkfzzu/0flBdJfNry
5sNoF36EV3rfLFDSRx+FcAtWGnhtt27jJenAafOljbTf8YzhOu1wgGuW1AtW8xftM4WswmHULD4T
Rxk/BeJJg2l8IqdEQ0/4pWItMuLW8+kJLeg+yxS4fga4lK6xFpRRcz0hwAlq+MIO2N/R0G4C7cnt
b/+BLPaVnzpcipB8fw0wtW42hQCbM9GPrY6D/RYQgXXWZWuhulbv+7ggSeXIYNzQDn+dYbFz53OE
rWD/ztHXK9d6QIC7KvEmgyb6SZcxtwWNhEFa14LFJNFzVfEgo/mcqFI/Q+Yv0BQhIfq1xX2yWFHS
1X0PjFAE9Q32k8mjHaUhFBnLGP+fzPm1oT0l1hrounKE+6uSo/EIKBq65CWKdr9V1nlmJdveN5Lj
1EX4uAe+/lS8KBBZL29ILzkAf1REA4S6lLo2kMTdYulw9CJsNfwzawgMBkALXNl4cyyTUXSs7xQv
yXXc5DHn+Z3vWxoyXYxo7xPynY3SDN4LHCVE7jeKZYydDL2TTE7bs3OZaG6VBM8Ss8saw04t8MQr
Z2zavs7mDDsQ5dcQP1TNWj5Ob5BqAEqcMTgCpXv0PYfiRIpNJFnBFhzYvnEZxhNV1wV76p6SEcR4
m3pNFr1Kfd8XmMPrOoy2NZhOpPNoSOy3WgWs11QYEAgT8+5oOy5OaXx3qbwINXfksOy5dM4gH1TN
j6Vfye5d7fIoso3JrXAPbqKP62Ckmioc462v0j2bgjB/8ha0RSupcHalyfMCePxFJ9fPYKp85NGe
p/zEh+4rTnUgPuF+HiF30FRCHuT6FQF8znbhLcFQG/EOcGrKT2aTlwZG9m7k+9ZLQFNpzNR4AnrQ
3nBWj97vlMvNLfBM4ImcVTEUhZQidl2cBz3JwjInz9z40Ghd2B+GtdllAYy8miSYpJ5C7ddYEl0x
ry5A5qVqDCMlDMhXZppMnlS8GV4+swO9AQHO/MhkjYhZK0pDOyN3i4OavZmIeKnBv2Up2AzYgm+Z
JAeAPDbTbwpPWp2Zab+e9rqsVFxgRaNTZIFG/HmgkmsE0hsQqeeHEdkAx6Brz5+w6cyervFiJzSx
Sc2Ji5wNEHXPoOBP2weMdYZill+3qdzQobYRHWEY/sbmPtjHGNsKY+ZTWMR0puRj8P3164VnlJJg
e5uMWgls4iZcWcxlzpiGP1nDQ6PkqJ3nJCDTTBhrWCi0L/0jJw1yiRCPXbYZCZqf545Zf4bmVWlg
F1xyXs1kuIq+JoquWBOUPoy+AHWbwGwOjo1lm1YUibLm5zNVpUmKhRlmvJuirktbCMxHfgC1jT5/
yUHD3xUJI6DjlbwEy1K6czZUYw8LbDneWu3KrQ6/0atbJV6XgTzwUHMmAcx3/qLTOjM2gh7IX34d
NYSVJYFwRvT9ZJsBHMJHNF1N1kxZouxTP3hV3oayMOjy4Rpo+WrCchH4HNICqL4F/LwEz586Y4Gp
QEoyz8OXv2FmlJeLE5uIIWRpEFgH7j6UB7/qjRR/7SYEJwLv7PqUmBd/d3Vt9O1A6pvepUVt0J6A
RH76hvEOmoBK7WBE3KgEgQV+/j2wnkpWDyuCS6fmEOwama1FcyvgKYPS3nzbklWdMWSDEl6NnpC6
q8M8PMXVB8jkPpHI2UGWUEo0H7LzeDIFbWEEKVFI4YVZ9YhjqXBkH091X0zjKIrOxKx6mKeLbRJB
dpDHpvlACM0X2v2Cmw/wP10f9ZqG9GNX5VJe3ScRZUJa9uEDkzVKcbneFkWRQJManzTRtYRP0mM5
05El+/cs6JQ215Pz4RLD8G0hnov3Mb9P9+/sRNVD1QS8evjW2qspJr2ZaYe6VvD9j/UC5Fe10yX4
sWFTKV3IEb0Ars0iltGOxRKPUyxU3ydezeOjiUorBbvWW7tuNoSX3Fpo8OUDRUjHBkZIGKPW8BZ4
hXj2zHqfB0ihYI+DqFpQYUE9T+YufvtqGkZAzET81F0NFR4DaL+yDFCTG4RAEOVhnKc8nTxoXaBN
4zU236lKcUjrcf2Fry5XeFpLkDX+hwb7ykpbNcsWHQtEsKhrMiE/JUPHYsQ8BI9+5jBCcjoUfM2k
VObusz1dX4wKAM7Y5hHG9PDH3EoSRl1J6yMzxSOx2V/E6IxXe7FANtUGiJRETq2EuQPy2CXBxdg9
3nVwHpdlZkdgSz8TvYCoC0zX7dUKN0S5nebJyJ23VQkPejylzKWWxjzmb0T6HhceueWJO9bWOZqk
+bXn9ncNEY6QB7gEf9UwyXNOeYXAALmyvJhzv6vDWdpvWUz1Y7gGJm23MPOTc6Z7WEDldNxjXvaK
mdU7uZMvnXNhWWlPUF1hfKMdRBQEFaxfC+61h5ImMdhQPFNNPtBqt3ZwU8LtAy3HdYx4djqj1EP4
u7cTUcvwfAe44K/kRTZfubySBqKMg1SmGfioYRJP510AAd8zhWX+KQXGRBkv6VJRx8UeMBMUa2KT
PtjpnUbKtxPSssdxJjale07GnGxyLieOkeprgeeeVxWKMXDVTYH1iWUNKpsD/aSDC1x6aKJyZPSg
sLK9t0++NEf3tITZy/kaqVZyfcGH4AjnWp97BrqBCQE4N8JUvec1vIQA84uKgQgO5Eze1TGUxu/e
27/51srGU/tYW/rGmq2jCohukqojqeTsf6/bf6nUsvCGOljjzhugISzTCDleVwBj4OyYw8RVhXpd
3Z2mymYWnWKBDsXCHjS5BpK1NsxjzT99o6ikneedop8eHvQzSPHJF+Wz3B8XfLTtKWKxrjgYB/i0
hmN69SteZoF1r6aVSgYS8tsNc9Lzuy6TQHPevEhwBx854YzWd+yWAshg5gkT6you2T4KmZn8gJiU
SZTe5Qz70P8zrDKN/Mz+pFaIii6xsCD4waOJsiQLuvwfl5tbI/jgpo32g/gZodQv7/sVd4FY6I/L
mA9WIYbAW/f9BcAlvTVc0L2/APX4CC4P8N+gkFKdpOVOQ66Iod8nDeXJ0p/zB/Xp0J+/Pcdfj43Z
9RtQGVNfovDQhZuK06WJm60Jx2a3AX5up8DUYIHFmbgP1e6nO38DLvdp1Nf8d/OncY/dSm9M/u1x
BYfYq/7Mk6Q0y4nX1xegqD2knYBU4mPCJiM6fzURwKpB3Og1+vkYUFSBr7VYuNqNo+CqAzYSWWN0
XfaPRTQOscAGYq6pbNp9iZI6R39IFiS1q2HMey0QjGdaDlgtcUT35Bq7EvEkPRbrKpA7bzr0HcOH
jbj+as2aJV1GcIumVUfV4ERKRCszGdCOPCB+FTtYMr5n2/hUbE7zH4y9WC2MNL38ckcivhXELp7e
YH8o9ljYd0uozx6GvYdhu667AVJuozMkHC4M9lmEZG4Qqi2ciEMuZL0DzQe9WDXmTUGrGRlmbu5Q
jmjSEN/FEl2F69yF6SovaiNNaO0hZtsXFzVJVSK2kJ5YQfmdYD241QK215OrpqqM52CqXKda65SQ
2etehyqgVVx3BPUaMI+sMPPrQGXjPXpBmAmj5otbwXjOInoUxU1x4ZWjYHcLRsyRFuiwXsB4b8o6
NiQ9uHmtrzcdmBOXyQZPOBJgwEV8y0lwVE4zNyblBN3FO5Cz7MslX77+izAr+pU/9XyXAeF6TqPH
TwQbr5a+9HMHD8c8DVN0TsWV9nhKEH5QOEk/kzkveOqdhXSapTNW31Z8iDAFYAKh3cinqttXK3Xz
dft2QjJGck3JYW+n9tU032VZY6VM4+Ej5gZY38SRw9PvyqP0CC2633KFDdmlOaTkk6kM8LzLdeMh
9UlzJW0vNehPCd9pZCTCGikuVH5vB7yqwGzPZsze/5HzyA++xzurXgKfRy3RtJuH4dvhQ4ecTQrg
bb+zzG1PU+RfWkNeK78aXFtmq3Xcc9PFIJgy89y90EiK2/wnZOPa5dZu/dSvGFRWsapA2+dEzZ0J
8dUHBdMNonoBKBRHqKKIiTUr4GM70prMx0KPrKtqrUmr/P0BLOve10CZrnpc75kG8nqIuUthQRSJ
+xydacrePLgBFWMAFzWPoIOfuwlB7uRpCqwLn1ilIAG8b4NpoN6C7xYr8VRbvyO7/dPoOCeSUrzO
h+ePcwXqa+J7z+xzWAA3bValn2FbNJFLLJ7uxJCtDzwQaV8Tfqan/3Fk7fu3lIGu4u3hFnfpiOaK
w/rMeGW1TM6fBWgGLwZjZ0c++ndxkC11b/Q+3ri3YzafUs293rtKTEObTrJ2AzrdfqyZuwS8a64f
VQ572HegeTak60Zlmg/iSHUGltAUrKSxMfo42Z4CWOjxZZYKbfiGPD4/MTeWHWwl8P51KgY2adhb
kC3pr7hY5h2ypM5MkAvss+TFf90w+uuSPiHwyvCCMxQ75WHArA7tIv2jrDUuUPWn29y+Fj+NnLTw
ZOxhvxpw2mBZU+5HnHmNpg0daPOEVWA9039djeUOqeU1QED/YSyFWMj6CG8SPD2jEgqb7B1Pmeik
i/1sgmgZ2F+r2h70T3fKPajDc4Duki51PUto0HkM7nxg/JUHsrBOtU0FcyF8GnTI7rCXg8iKr1g6
c+bEkDUeldPcn46mk4nIHNmgaCG4dEGAvBvTmDPWIVsNfOO5BbWcmLVFe1Bg3sEj8AHVLHkTKj9e
j+GpASMg1IPhLp5c24zE8u/wvEqLj0H5oBrg85HYpsBGkMNMrXPo7zomHP02eYvGezl3De4o8+4a
SSFFz2v7M5c8cFkyWPbGdoJWRcV3MEt9PzyWPwYk/yjHsNBJmsdnJgCVlak4aexj0JGodABBYHjh
p1w4gBx0TyLreaz09tFXdsGxLSX+KCMcP/OFDIOfUdXmKN9+5pqFHK5VoOTKUYfNZwKSAPWh3V/8
LokcVmOzGQEGjHbcS0PnvJOvFrfPj0I5gvdBi5NlqeaueW7REAPu+3VP+0othBsOAhet2JTiDhc/
JctO02as0qRW/zb4caoZSPElRhFRwe/cJY1N+Ncq8MZs/C4Aoi+n+FfHQPpUV2trx/nAleJHGkTS
6yJao7jnEij660gyUvvm0xYKSzYnCxmhnTKOBwqfDw2JCjvIEvNcQF7RpG0Rbsw9fypszHaKn78x
QQj138/b+jCLAae6K7wRCdRvXNa7mx8CoPdcGrnUVYF1PKaAgJ3bnirlBn/rt3jmhxciKdsLNSge
a1uqpSbbWfWnSOb/ijHYkdePaWTF5EjjFbPadQA3fbjEI5BHJzQDSkKsxEZB6mx3ccR1/WvzHLz5
kOXpdX0AyaohBPlHspgWMUGcy22qiWWyNuzkGHRxsa9W2Gm3pdRUpY4aKg5rgsiB5rNagyVCiLYe
Z88RoZapC78FVYvFCj7GhPqkul9s3iRtkbUcR60bhqGZotn1zILa4Y+kgHkytDj8RsEfs+NDGHz3
BhZ8cWdvSFRiqliiIJHHL3KsFOeZcgw80vFeM1O0pxlOHVPCSAq/siApP1dp7YqFeYuhb6ha6W5N
nBLH2I3GRi29fPzPyZ1WvLL6stuqCbWtJcwiKRS2wzJfBquSs99FtRh9wTiT80faOIxL9igSvR+D
PHA5wjIwWJwyD30JF2xP/LrLZL5UOe3pke1Tiv+YDow6QuP1USfm9R1sQTp59x/2pCNEjlNZJV+d
cTPI4tixfMhkzc+QFsmEQBdzNH45aO7dxWeatKrpDhXhrZ+q9mOIHFIzAbKbsR35IUGeulBmICth
uEzAIzCV9VHnZrO0YNjk8LSuiCbxumqQcStKDhB10JQ5Rs4ICTAKcjhcq95g2bPEv5ESGKRysasL
zhAYEH/BzGkDU7Izgr7C1BZUe2AAZBn+U/1hKgEwPHM9wCh1XnIn1Bs4KNxfbjPv8DX3IfroBEv2
Fjnp4qIamJLu5SpgmrNaeQVxKPdSeJQJGsd94mzFEu1ChHfwyPJ91wOvXsm+u8PePzLueyCpGPJ+
geQrjDvXQA7CJDJgrP5od/iFPGdHrwOd26caAYN6o3/TZXGEb8Uc0BIAmVvzkgFMnM12jXV3++lP
wNnYUYakoapWSlJAKkJGedQZLLN86gbQ8pRSj9lphNWaofe7a/WLqYLIhEY4a+Vb59xTKmStg6Bk
+dOUOaHL10hBFiSzH2utDk8CA39co81QJEcnYSXrknHIDUss7Hx3BHTpz2EIHkvnQkzO74+rGkKW
VZncc6M6a/ZjTaoBmrNykvuGU+ZVmoi5q5bMijGQWB2vMeE5PS/OdpWqGH2CBwz2ZefCWdBkMXSB
mKxrdC+eAKdI6r9rDH5yFBm7lyW5VBjxhEPnDPBBP5WqVKiNyYbe4rwIH74BqV+zQVcTL2PwE+jG
9oZfZHjOlhVNQLfBdo/mKD4HO6sF1y5a7Kv8PY+FjWrEFfiWp3aW0mSE1Ms5189CMUgxtDa8JrMo
9/xz7SWtFbjqurUVSk3GLi53EHaBJntuYfyD06EcUaYqMBny/wr6eh4SEM7f7287OTkg987qjyDD
kWlWHFyzN3RC2cP/ntmGIvq0Go3IEmepp0gLl2IT43S35zBubEDvP+1P4vIvMGPGqbT0sAc9NXD2
t6FQrgCXokCTGO/vm4CtN7c4BEDf1qSu2nMeteVHuTQ2pkUZYZqhpdBpdX0dJCoyORe4/p3SlYQX
aEX8FAuNZCOeBwHIpx6sGB4KPX2PFHNQB7zsmD83qVOWBB7NQd3vqsi5HExD078CBJgbCMr2bzEr
G/NRmVow9Rd/oiyRm47Vf2uAAlgqLVLzN82pe6utVhpQh065+PcdypDYJhK1bNnvK1bzAxWsguu6
jSEy+kL7z+cSGSeixyy4EZ1nmJUmoztSlekuNnuHa+auU4pyWnpXCm3avYkFITNCiA/zFIDgxWyX
C/XyHtWVYiol2w7rosXMO2x97sruaQjlKS69eiKxGYpMRh6lC1qET2au95sacCBjsnicafba4Qvv
6VLt5+fus+DygYhTce1/fLXim1RfrQCIoe1GrSZ7sc6GEe+5oNx81AvEfizUMJmNSqnv07slN7DL
POtPEyvIDVx8ZQL+S77h0fAzasWZk0bvJYS1AvIJDkA3SoKUVBupQULNzOe1KO1nOXa6RNBaWW7x
yoXa6c9F2dakiE3wTuBBNKN6Y2e4IYW45zFoLDgxiLQxGlozo/fXS68koNtb6Llq5JuGkSmmWs/j
Sbw1FAkl+qK+TvDEt4ZkmUTRtsaKf66RwZmCVU+MtPGCZ1djW7OPgXOUhQS+c5l184B/I6mr26Em
31Aq2+V3Q/uoz0ZqTgrV2qbXA8Udk7CrwEsYldZlYiL92c6BlSHCtP8qOf0LDYYeNKSY+naq2aVa
Uy021APXzB6LCtVfYgV78P5ygnIdJWR82B46UBx03pmgTRihisRSZ5cmOxN4kHqPFGeuRXVeWKcv
qmjYrnm02esnaff2wS+3LGstYzxOaSyYMVdlCLj7Ur9wpP/qghUTUaBMUFbMMPSByy7dIbtgFJJT
TbEsZhUbj70aDUJekkmuD7Nm3a9KMBhPhZIXsxRR4GiTpd0r6JYnLbfvMrJ255ZUWPCBPgxMy4g3
22rMFa/Oq+zuOcLy+eorS34Jr8UpJ7QabwrHo3qMRawhq5EJ7WX3MRPQi/mIxZCNSBf053zBDFCB
cw5iiEmu85EX6+uH+7vip01u3VPHFCd8ERDQ/cxSlvheLbeb0BuYNbVwBuWB2+bJjSU1iqDlNJyJ
BE9DcZjxq6wnYkUrsemWvBRMbNblWOPT6YTmkc0MzVrWmeKCNiZNjl3Ga3i7jFsqkinS24yQxosS
ses9kizXEqnUA95QZJg3N56NRNhBIStuw1XQdZL1v5f06J4XWh9l57ZacvAGxeFbH/OQ1493mZ7s
kZchHqgimYN7WAoz5BvMSq3Oozz62fQ4oqBplK+V9+GXlsLRdQ8fzLOGKMtR6Z318wI5ApodJA53
q0tjzZY86+LuO1hXx2rL1svciORBkTSgTj0Okjksy2cVem9+DZbE3T5tqOXtM/xNq0LT3wnN72Yh
eK2GGiFN1X8aWkc8kaXQ+vcWXTauPBr/hsInPqM5Yzajogq9AR109nConINiFlJcGK++D/Na4gmg
61w7YwjIe0p9vO0AisZUvkr00Pcj8zMTcAQUOxv7hdIMH6HFBBiCALYAEx29Z/y+5oAydR7iu+sd
/LhWQLv6H4HaYVyrmtv9MCUhK18GHdTqXXF5vlYyW5gnPkKQUU2Bcv2bKHhb33sJpnNjB7UqhdHb
OFk6gU3o6vc0PqKfzCJHHHccDCiqV7DoNLb62+RSNrbzJL5mNcprquKF8NYULgCQA6abkKak7i0l
2OjQl14Lo6Jz/CJmNnlT2CoNGkjo9PGOQvlND1bfMRVV94DMUgmZ0swqYRGl/cSQ7pdTijsNVQw7
Mrv1YLU2hCDRXjDZH+c3huLOtgxXK+ifn3QtQHcZQa++QrfxgBolO6AfWuNrvfDkAYE0pfzRHBWo
OjxkorXN6eCD4TgsiQZDwcnsmNfVZfxMje8yoj+uFUEt1yF0Wwhb0YDIRRyJVCzXy5XTMn0NWd2N
85+BDlEUwq/6BUJbxMcdszCkpbVwwcWm27dJC/nRXUXZnLZJH9U4ALvRxcLDhYuDqJQF3E/d8hdU
CnWgGp+o1KtEN4HKrJ8JgOr+SjoJ0t3bU9E4ACRexqo3nwqCIEO9vrA/RPFA3GARSbf54cIeUaCd
UqGZ0ipgaiSazRdVHFcXR9vklU5zJhctwwRs7R3VR5gi8Oy0zUuvggB/wmfp7VwfUgpdaQxCkmME
wtueEPyhGafYPZ904nbI4ro+PVYmCaBGu8K7Ec3cloxSuJQcI6sRLo+u6oCDKqs33uWFgr3GU64z
Van1r4BRywmC/vZZ7dv+UHAfZX1P+JwYXPK6+XIG2ceT0tNV8JgOafJ/WYSE8wx645tRklEMRKAL
BYggulktJHzevzlJOd8VZQCTy3jQRz8P+aC7AVXjGyz8NLrPzrQSZnGDk9GlFaCjT/BNEAK/Yodn
74TA47wOLImjtPHLJ32Tj9qEBHz+gixBqZunDf6195yu/dHUa3bWZs/+lGfS8+RaQxl2FoECXfUT
QMWuZzQdmfmXGpA24aJYuIoaT7vsaTfAEtz7j1G0h0N5c1FMMBDPiog5+QjKoLa3aXkfABeiJpLf
T+DdMYdFWUI4VDmBnb4tBYxzzFCXZIuOdyE6ybi2H9XlU7cN+f6nVvtH7rFqRuhwvBRf94lKt7AL
/Gl4p3l2EDmHI1iEXCA8zvH/bW3YUHiuYR6FTcvfCQwjF+TuKojOYOXAUUvDO+A3g5T3csoZYJti
W/4Cw+t47EyHw8eWpPKvUuphzxdTWOHRLE8K3uMQoPyrgcb/H9WtvpyJXz9bO/PYNonCnxVUuame
oi4FDDAOzn6vsZTpRM2qUAWwIuvR5FT6FfQqQu33mEyPCB5tiANn1e9yRbRQR7WSeH1QHcSUg+cc
usKmDCt2Ug5CvycVuWuMT9SuVYLzLDUbjdsNIfhN5GDeJoJTuH9dhuC2ysVbN3SaqZPPx0IFCxYP
nRuXDLB/vmfhh30/remz1in4staEQwY6uN43fki8ozdY2jp9wgCdp7qse/n/xwnYTUCbJiqbZiWt
4A+x93lK7rdSaRKegQjggXhLB99YX++15QPyjdoRmmLRRWgi3fIEWUz2uubSQNCkQ43dINX5qPdU
Mu+m+x9uAaNX4WQ3Xl9RHX8NeBu/cmWOjTUxIuVboDw2V07vAvWu0yRamr8TfXLjCFvK2riK87du
ZxsxEyrbpUekBuN/JbrSZjCVl/gXmtoVsTUJC0yJJK7koX1Kfqtort0rkkVtnHrJAYy1q5tJT3m5
F2Nvz4fKRAxR7dDfuWR4h/ZFzZd+VvvfwgKK6VCYHlE/4qljoX4KYwy3yTAyom4b/FwFxPCwrG/s
AgpGurp6VZwJEVwkU4t3FfWHVN9NyEn0TnQC7QDcodHckKcNF6Ij2i9zKyixNp0JyQHDwM8BxZzm
yp0PGOtneebMB/pARTj7HhaZneC+bO3p5ZRYemGVA0HBpXbiZOoi1sG7EWJl9EwSWX82fP5ccf6D
eeJzcz8SX0P4CF9HKmEEtAGzqoDXO+SgobLrFEk4euU8lcLwBHJfXKAHPyEDP99veagmLeA2QZRM
//imybnD/UzTL5xcGjSKsrhEalWm2BxRqqZhFVaagECg3Tt1dqcV8V01FjJwWH/g9KkRkpxYS2vC
O4t9uPTeHI+qCGtPtr0YTS12JHc3+TV0uR7gs8GnXZNugIXyGAh+/KhYw7YJND4troxcdaEwWKOB
cPiqJ7F7cfZH5Ia9/c/bfiKHjNA64wqGN2Vu9j5rM0PUghuV+81VT5vFfDYFvU/vYe1Nuw9OxlQg
By+pGAxGBgC8qjTl7M6jat/fSy7uUZwX1/+Yibi1NZAAN2oVibNL9K6DMxBYNrbl22RznZFvgTqj
2VxQAjOmJNhY+iiBaWJ595f1XK10kFEVVdFr54mA/HLQE3zHjrHpX4T2aEc0AQ83jmJpD++fxVtA
NKoFhi0ssfITaUlVZAtkhedXVzUzTetaKFfZfoR4byWcabbnw+gKcOYhXgehLSFfIed9kRj6c0iG
40/PfwQ7XDLuiM5+u40XH5fNiO6IdsQNyPlT4t7q4Q0ucl4AWSXvNn9zvS5LpZA3HUehQpu9APbJ
6gnJjD7WiiHDvoGazqMlvpzu2Ntv5hW/Mz11+RtAc8FUxCvAr6XowNv0YMjOTa8KnxVqLEk1XesI
Fc3YT4SQdD6FR5Ib8QIjEpQv6LtNXto3lmozEALJJS8nQLa2cynI7wpzAz06F2nTx+fUtWj0gLRr
XdEy5kpDMn4/YHmVxbbwathUYSQCuPYbdQZRpTbmmkKH9l+a+NVUocURxTaPBnCV292d7DqcWyhd
daHfN3TdEMrn8EP3JsGDZf6UiKM4SlZ+nyB/Lyah+XWOV+RJHX3U9yXL0+iiRk2XKurHlL+ok352
O6N00oEDNkg5IrpJP1CUbQ9DLQvlE1hR1XtJpxfj6+uC7K0FufrniMPOQpIRp+lszxVDT7Mnr+HN
iPJ45uX2j2SPRxhw7wSQ6kMkK1PzUCiduxX+lk5jFgfuAfW6i4RF/Se4O00MP8mytHdd2QggvOVA
LT1EUeRoiRGVKMnd0hU5vWIOXVqgexeQJHCasfywoja1VwkaWaXi7bdw5ubqMTidzFTTA3byBhlh
ybq5PsmEEvnAo4YEIE9ZhQu7bQVAUQlFs1iyUZPvn6jLSjCPdwGe7igQxxM6I1QJWlJY4rZ9Jhgb
1o2AJAMeNVoMkMEutz1b3agDLXBnV5VnZ6ev6n25DOeTvQhot2W060DdO9bnZvEJgI9TH/nffdjw
T9km3FOFSQj7qS3jPNZ8NgdyJ0AM8zDVlqgpfBsmmS64M+GzwuZX3jQQ7xYZvl0JM9SEBUD4ORqt
8/pDzqOV5XeT52rmkHjEyb/mWTWl2LwEN2a8Q1q1Qn/f1vEPWKjLe2RX/xQb1/uvaecEpy1NXZn2
kO0F4cvoCmnT1kApiS7O4F0gC46qded7w5rV3NAA0AgVYhCcnz6tNex9GWwQZB6/k12Q28TUwOsJ
amSPfvcqpoprTZ3e5pc4hSGzBAMvELUuIAlNQPbPKmVAjSpdalH5L0Ck7P5sbU0fNKsg5aTc7XLX
Z2pYalFuM4G6cCaqMaDehkmFniT8MZFybdV2PigM153TocNKSE0r4qYqlbjB7zY/p2HC/aVi07K0
HKxNoJHfD8SWEzllcpHlYHRT4g8lsWkkHiKeQBhlU0PAaY74h8Yq0E1kXLAwu7kHdftVXCBbXS/E
fSGuKfUtIZU3LfWY5I2cTQWO9XiCuQKkpxmrK9hrSmZkIb1dNjmwsxnfsCRRwuGH95OL+ubnvrS+
W/ws6ktTJJNBhYBhLMIo6fWNMWw+5KpDwLgIf6ug3e1WWii/YKx2vpM3/7Vaq2U26jLEmF37shVu
WT0J1OT7w3BJ4USKh9ZwblQ3D3baxUnMqh0yWEhKzYqrdvB06XljEe77N58/jNtHHp0auZJ6Q+lL
wBuM+9GPQfe+yJI6/3anv0nksRwUkc/uXw2+rsxZ6MDngzeiT/V3ztibje3Nn32wjSY0OJ6mTYD8
zYOVBF365F5nCXjwMMZhvqLbg1XkkRvKHSjL3nPzKxr4x+cLzpohI2AAhCXJCqzc0zDgsYhr+kqb
g45tBXQNIAVwLaxU/NKFEagolwP+yE2QAN7nqLsRXcnjTKYclW0C3YASDB361aeX4DuuJt4gob2A
0/uxMOLXULjjyG/KX2iVVX7da4K/XeJ9zDVYfUl9Nk0tM7y9lXhaxoeDQ8KfYxKzDPbXkdwpi7Yb
K6m6pls/1joth4U0iuDJa01+0cU1eXRHFBkx02DMa0dPN1F6a6rhP2diR9FQIuP2fo5WqRhwxVDA
TUyvVsZn5RE3OiQSEvQRQEIT3nvOsAJ2hjpdGaHyG7zhp0/PcPSjuKWTfpOBgSTyeJbhVcYEDNTI
shrYR1afY+W5XR9YuJqqsqoZEbKlzyHnP9W3oSL5s1qVv7PBvZdLL/FlYro4el3OsKv7bNtjGSR4
nDOtVzIsn8bF9sYUrGVS3YI7QYy2GgXHZYBMuaOwJlXCS2H2LWLHP8ffgxM0PRwy3F6n3LbAuDTr
8jUMX870Kw9fqZvRKTcOEZWtyeEl0q90NB3FeqbGSdeu3vCrUFGP7sNY4INydqO/fjIwbkYVbVA1
oHDCZqxabQ+ZqbsrlqsssP9D1oph82msNScybRrTrMj2/3SBphM/+DA58Pxj5ZtwhBfFiaXmCs0a
oMD5WDEq8Fm0F2CXZDwnpZaJotHx+sSwHN0iNd/Mepp7ByXtiXDyRhZt6WDe3sKZOgjo/IVzFPi5
lzy3gHz4ngCJz8jKGpfKZ91nYApQq/3Ml97iTuSl0enZOjf+4YNYtSv48EhI9JzBfagOSeStlcxl
PuSobTw4SKLwC1vyLAQfHlY4MYY+YWrcvnE5M9H8I5cVfcL8uK5v2vuqzqS6fddUOYtamgdq2UZm
JTsk2vzNLugc18cV2s9yEFXNXPXbq7WJFauvuxU9YcST2rBB1qFiOeD0TeWTLQjVGKiTgAF3hPEc
PIOHKSa2mNi8l8f9qO1zw+wGpVPaLquRMJkKnuJduzfu0llS8mAeurTiINNsLFyR+/IAJaROg/fg
hp2RfboRbPUH8vB42DC+MvrxbRg6mnk/Fr8g+NSVOxETzJMqNZ9PcjPDPc+av0LZpk3iyvXpYF9l
gbvXKHax78CQ6gKI4CgfLGJ98g0pxYSvzP8knGKiojWmh5w2SEjM7ynohl5xmRdvkjoR9ZmwULHS
0/ijWy5xmN5jGrGh5Lcb1MEcbE+7bCBd7hVasVnLNaUhGw4wu+yfdZgJz3KD2loG1wR5NkZnYclw
yT4JeDRsVP2W21aG9/wcSGJUcNWf6+hjSRwS67dDPbc0uYu/ZEpJb5Cf/bjBiUOoBNfO7nlJ68Am
EJ2cKCX0UgdqZ8wrOPz3EmSJpZzveSPpb5I6f73WvRDdzdjKSxJdfaPofrCxPiam3ImycJzzYrLj
Fojyj+rjwx8drnGafsL3iLswJbbR2znSQGAbEIXp93gveHrYpUixSialhUe4hiUELO3KGVw7+DSo
qCsG9Fcqzs7aPnMV70rIevhswuJddkJ6Wl2taJp/KUBg8xO25N5121yNsaxVltjb3qv2iFsfXkJ/
jB/Z+Ty0hL0wNczQMrVRDTe8DmGEMuH8THPLYgiEZR3qqAv5wYM5Lww3vseBV78XmRpEfLcd05wu
nyY72vFC3QSD8fc4pTFYAnqi0rqemADttGF63s2Ks6/FoQd17U/wsd24pQcIT96dOA9YQ3Tfm7Z1
QsqZIjQUhwtbOe11F/lNqrXe5yvDt/tdEx73GCJFhwJfdz4j2ErZUKVduRfdjT0wZ3cTpwTe5gbP
h/uuTzRMyutIUZrKSQd9DnJVIlogWX2HFaYZk9DCItF/Es+M9XOqTvOks9RJY0AVK4wW+us66n0m
xdzATJu9b0jnICgQtQiIf4mLlPLdKYSDh4gUyOxhqGcVSaS3zREFzaTGrPW9nGDrarmO2SzDss2M
HE/Ro1eqbsBFfmCgIeXXQLpHVsK368j+5DBwh6rjUaKEm/mR0OR43L2ClQXjTS8WoGWJSToYaJKJ
fzu2xH6FFPMaHrs3lnUi+VBgxbgPCHx5iIYkQRE/HwTMcJlRmVV7eGDxAgZ0adMyMtlAtPgs1ptF
nRHj0Lf5f8JIX1VsGH1KRISQCPq2MuGBJaL5J4U/KHlB4ABxuqqNNgfWKiXwdqpTRWMsKosnTfuo
9b0xR5n1daQuoUiQUa6jH8Hj7Er/FiiDm6IZe1cXkMBk9vs3/KoZPVc7LeqayZSIh12AR/NkwSRB
xNxECWVapD3gGvzDU8ZFGv4z4AyhBg+8L0Bj6UIlHSdk+DeY7bkv7nFp2WkkLyq58P5adD++Fq0W
dIMK6PhlYyv1mETVQs5N+5WtXVmX32XB5dAbI1jYhVFN0uCd5Q/dreCyV7FlUhcLavGm5GZz0zIq
gt+KAvG+tF8QSC+KFh4r1AgqSAoNLRl4aYb4mNCLR/Kf5RxRH8bncJgFwvGMfQU45Wc0MrgyoFv2
kEgKMvNJ4YZu7juHZv1NGbpllOmLoI5+phj8BlPrXhj3EmozEVOWJahSQ42SKLwsdem4N/Nl3eS2
cb4PU8+3lwaluMGfVb8+jx0HC+ChfeJ2nFcPMq+IDDzgkfzDe6gm4R300nCPtPq5MhcDcm98b9QH
CC5mWhd9m/5H/4thuCyD24Crcebv11wHH88ILu6NXTW0wSftMEPlSiLxluQJYu03nkmJ8gcHqhXb
/+JlauceX6cZZifoA3eOrlQ7pgbit8HSWuib9g5CpjY0eg7KTK5tpfeFGAETzco+CjMSrxklWtmY
wQibQ0WJGf8JqsTwMs+y41JHlvbd/fTl5C2r2klyzIO7csE7y6n+cpbQyMnRkodJHVftt3Yj9gGH
DFoC17mydxAsIhLb0Wl/tsF3hemh9xTM7UoGOukj3ib2F4yNi84Sb7jbYE+cj6LJOXuPRXYeZmnI
ThDlGJQL0UBLRQqbD+FCoZuhhVO5HcwxEqhwzjy0a8n+f5HU6sfA9iBcL3NVEAoczy+ZqrJ4hFj+
v+IRNSOPxqJEAwFs//UYf6vgK893MmeIjG76OopVIInLDcGLoNlyQyI6uXx+u9qG/0d0SitMRS5S
Jz0KW3ItLZrUpeuGc5zY2kd5Ye/QYmfLJ19AtKIBZ+JHQyM0mEgPLzzYaE9MFQFTT/Gs/QcB0twK
oUKGhmrmH5v42Rm5JNDSWKcBjz5w50gbGcyP67QQRmnSK6BtghDzztpv0CeGx5mzQjHCV8oqpwqc
3BBregXT+jY+OGwKTkJPYi66qIvXDGpYJgtllJy5aNB4sDoQy2PCtG5wZfwBXYhweLjj4WooVEtx
ThbTMLZKGZkdFSGDA+01Pqug1qGiPchsVS8kbzvSr4esJRherZpAms8kO+6cIise1ToMiyGxOgZ8
ywETACctR6lACwU8DO5fczb4lBKSDnJUQZYR/pVJPvg3VKiwNs0npovoYO1+STLFQt1yrP99/sGB
Th8ayHxrWksrissG3wQbwkI93wdi4FbtlHaLG5giL60o3Z0Pk7B3pJcv8OQWTtEnkDb/N257zO14
krWiPkacdotz49jjbrSuCRkMsjJxKH35mAEqisSwRaqHKfGADhOu7k010WrP1bjQaR9X+08h3yPo
37qKQoB4tNOxmlIQBcHcFindJ+oufsJ/L/KralMXevBphyrS6GRn7qxy85y+9AbliEwL6k8XDpwi
SptK6CMW3G3WpLiidXvDpikasCBPyvVnvmKnYCFajNLU0IvZlO4tIxX8XWXOyuCbtX1BbxmHqNuv
/zQLUKae8+8sOQ7uLqnAxjfBrw5x2ZPzjTL3a9Z19g8Tk13lvwKNX2rR+issLibkBR/0e/1mUvpx
aObqofLIwf8Qyy0+cw53IqQi2SAUZxuGr97O6G6LuQKfWBqMgBS3rpwEi/Lfsun6T9BLJpb0I+2m
LlP8YxgrLEZV8akzv8+LntgcQHwg9RCOdWH2/Fbf1/6NUheuCOQR2UJ5xIMnuWnJJeC2J4jotOJF
vBBSk4xfc4rDkEybMqBMW1Yy6lMLXrJzB1JoenkLUlA0wtGCbTzz4eAAqNoa+XmX8Ys0FO0Gd1Ij
OvtFlTjAvq6wxBq85EwDT9U/8yn+Amfp8lh42y48cgsR1A4vLnDUjwBH+Vh0eM76kFIVF8vZTtcJ
uBXAz9uALaRyiJcEP4AaeV0DX0567uz3vJyaZIXjxrWLe0Zn5R4HgPro4elYQbIgqAZhTa1x1PiE
vd1nroyTFvNfx8KMoCbiUwE6WeO7MB6+nXqNeujsCk4vyEHPnZ6lWY96bhoBzn5SIxsbBr1ON/8t
nuZjRZpsG1m5v7oKudd2MOYDMzfyzAz+cJGPxOucHgiym3OaCaMBpQSqbi1MQwDeuVNanWvmpC0q
FEQypqBg1Z0tGZx/1NLFYCvu9s0M/W2ceXCvUJGxNHC19oLlnoIKIWASscVyDvDq8M3B5HY1PxBX
X6ksjj1dHfDiPaebiUQ66JIOSMvhpKFaVIV7CFh9/7J+3Lpiffug/2bEVv1zCmd1Blu+Kb8zQnW/
sO3iLboFLOmfFipUOqMbB5iDd+kP4gNsAfwwzQsb3/flA2Qhi1mDupj3ZHRDCtiuZAoUdIX3B/wz
SJ+UjoMdnn/QJo1GvsN6k+Iqmd34g2QGVKTZ448SFKhQRxYJ4KNxCHsc9Tk0PNxq8R0pU0MV+S7c
eqR+fDF9XCyklKo0jKaB0LFdTn3q31fmpzmkowZCDAEQ4MnaKj5/RWi+TPSsvZkcRXYB1c6JBvwY
wpgPo4zxsMTy0qLlC2fpmtMLO2Ob45kOX2jk0nB2NKd0hy0DzfwaimqoRw/LhtnvzSYGMAQsjsVF
oblvRziqM/8enP5847JHM01ly1DWxv5iW57qt0KQhbPVVNQttzeddhcp8gumQYyeBft8B03JpDLf
UcT/cxfxFeZyyygI5nE7QUk7M17Ek73QbjZ73LwRGrjjyPBLECoyMwSudHPtvlzFir/cTg6MZ3Rr
3gXfZzQ6WD/kqAqQtqpGHKfG22FWQDMnBtYvJqMk63zvhx7IKMjO+7cQPVvDLZGwr1CEJ1YYcs/1
LPeQMKr0GH7c1WQQnZ8vJ5WoYNX0mhpfjhjL7dwgsgwtNLiKaSGz3EdUNF4TMYKbxDlIz+wgyjGY
jMlQjTDN2ov7GMUNLUvjahl/+vAQnNw1wBubwUpKJ9CfCvMbT37wqebeY+TrT3p5wciU65zsq1LY
wARPS6l+gRFuVVfsd4o59Hpap9ScRAKtX8gDd+nE/8Z3zLvf1gBqZEU8f7iDjQhNPsVFyjwqlNwO
MWAh1dsVRKWwYQanO/3+Cte/AEbygTyLJOe9dOM9rNdcTxIZPsKy9EYTdzqzOQNP4FFSgUSxC321
0XqB/l2vPRMZiI7ZANWl+kdqG20TzcmQT0pRcXPndsTKDlE7bWut4MZeFjC9jckufyhRZQTYPWyi
81i39cxrOAEjtGaAMMkYT1a9awp+zksUnKAxGSvb0ak+JsyLnpy5+llRNiZxA4lv+oSpdo5ZZ3vs
/KFsMJB9vxmefr2XtzmYULR6T+DfSjVUH5vsKMqS55yWPzEmgkY5UMkRGE5WYuGxuwtXpK+6A386
YBi8itMuRP9tD63O05UUF6Mk+obvuPf+B0ngvz/WFbxVw9dyBW/tOO/QnkVs/qN4I9MlUhM7lU6M
C3w6doidnFvjmmU6qEJSAsc2Mg/Lba/1P2b7bQQYW4kebeNpXBnNMmQjKoHKGtdV7QMf25lv2wfW
PHbZEKMKsH0Xhlcc/PFWTDlzqUPRKce0FM5fOneK90IFcWKrOjwEZZ+J2xz+fZtq+3HdVWXzg9Ek
7gXKHVZ/xuAMqSAxDQf3DcZxsQfUYTWr4osAQ6w5uyu1IRx5aOXzfe9Pg32XxjV5hnGqSaulrkCx
W/bQnXDNhzax9OvRX8pfvJZPbw+nyLrHMQJsAdo5yYhBDa5ja3OM1rsElYs0XiCwCmDTg9JbVxDY
lN+OOZL7k/trldVy9pAJssThNl5VW9IYue3uiysVk4zn5PBTK7hCKwyfI2v0xu/cw9PeSDULllXJ
2WiF2KtH4ACYqUfC3ba/6gzd+Bq6TI1a0laTVJJdw0qENhbblozdwYjQa922zwnCB9XWp/1GBlMU
fV5BD6u9h0HpEIHSQ1RC51+/nE2M38N/UeVX/A+FFmMGmezAD+m+XVsRYItwWjPVMFgqLcS/nE8G
/plit+YF+1NrzPeZHNYfEIZiP4RoMxIZ8odLCYDWTiLW2sOH6LIQiAiIhLp4f4Eu2T9gkSOIVu11
AVQvDsHOpffQAd+1pqDZMfVMOAGkmc1VhCgo4gwiZJJTIwGWOPzq/70vqNFNwem7ko1HwLTPFm09
PTSxE+/0Aa4cxA6Jfhv0vfDLA92t42Y5EfS+trakHKlJ1bM4qANs2ku1Y2onvZZuhmESxzvWgZ1O
6qoVvucegGh7sOrbiap6dWb5WlzdXO6eUFh7K9pzfhRnV8hT6Amo1cLzRe7YoCioHqezWE+G2z9R
i1hOBakJz4h08E42cj44bUdfnt/dBl+qm0pej2V4sUcE+wTvoHRZZs4kYbd29ABgNDWnUUsSfdaD
U5plOcUMPL3y75D4HTsx1DnE3lxEzrn13SvHATt4HVMrHtSpgKKBaGw3Q8Y5HIl++mXgyQYIpYNX
pxU14BiJFPkLFOPhGx6bWFADj6vChvlY64oEyJiKz/ALpHo4HKIRarEjlqEqx9/UM7dinuIf9//K
RMov5I1kLZ1dpgSMNRTofcezbWemWhwAyow4TddnE3suZ8UyG/zYHj0nE0BlmIuZZsSmdVSfZKFT
HREc4LdDInnIzrXTMxShb9sbMzmAnjNm6tdne0MRQvfWuQ2zJvJ6n53qQiWWi4HWq6QLOJ3spDDz
gGyumiC+QUvGhp/pEBPbIEeRiCMMFsS8WpBYFSZeo+MsQj2ZT1z6KIdBgqnhyV8qgqi+UL5DGWTL
BCrHQqesqS88ROXgYi8XCUhyAFlOTidaND9iEiOwEpdUz1HI+cXXEJNQVX/ileVB3tB2c7jVWrXZ
dduZQ+b47GNDEAedS+1GduAdCWsnTBOEpGMJ+Bd9Jbp0Jkk9xyOdHfNXJuanL+pFvtJjneNz0uvd
oeRr+AFsQybj/D/TIpVG8C+hOEEaI0yagohPN+jZE3MvDMeNLs9sFgaz9JJ4Qcdh6y2P2x6nFzKC
EFU2fXKbnzlfTc6wCJR8vELylnhKubkbTQD++2cHTeS3MMGx8DXBk61sayupBU2mpiiTlO5LcN9d
CoNKmA5JFEc1EsKX1Q4nfqYu7cAeGU88mvqaCcPcCjyK1jRC6LGL/sPVUe2yrYaWecLMfKjRUhMT
yp4kr47M2++R4sVGdcQuOPHvxcP2AJN1z8eTcjsUEfZAlS5VFVH1S0D9OMBTLoxDFfA91NDsA8Ts
gExtY1UEb3jFHyeP9OMhGZ+InWq/whikYj9ssl91XxnBXf4hDPef04r75aZg41C57FcFkY5UMKiY
0wYRZ2hotaUFN9q0tnfkfVV+5NTsTpCOcyRuBQcFQrcqHV2PyBlFSnwqgk39ADbQ/bxqR1g5lc+w
/xgZop7ZSrmqLq8tn8qDfSLO7dPd7Gftch+xc8eVu4ZAcN29PrAV3gr2ViOdNP3ziKdZH5hegiWn
4NyQNMXv0M5YkcXX7Zy5rPoLNkyqR664VUkPxdTNQOxeHfoCuJMgIH1xjpo0yXaxE8GvMSQRmXsP
CZdcQpte6LTaz9XQE09vsSac6uuyfZYl01yEMqiPs/wAdoj2xJX0OWvNT0onhM4hPNIVTu3EeKhx
EWGHHtlx/AT7mslbzH3Lziq2AEY2Dq6uIhDgghudnBnRkD1O0JjoIdmGJijuOkWIL3kFsCmvNzK7
ph1vB5syQnARLbLk1NKSw9sZLjHCT+R+JIGL+EFx6GOtYPD+XvXb77cfllxYVWPrPLNVcNUz3O2M
/+jRtRRGhY/OzUCHZ9R7y2IO94ZPd9DiAFsX+8j2zbtnvwpIDX0Z8sQCA1nLSNErCR9d6PmZ8Rue
imH03lfVWmX+1IwZpeFO4ogiclYnUk2aV9giUDfmfUe23w74y0GV7zDoMcEAIugDJTJYMJ5QIr3v
MJJ/NAHJQnYmTyCnSEGS4fYYbqApDGbrvW+rR7ns/U3FydIBmaMbo17nkVUk/KkS1fWXp4Ozjy9f
ObZtSKpbCWRKZS3Ig0GjXSNtOH32AequKu2YRmBjAUiKPEvnZSzTIzZal0iXOFZ50wmIyFIfCWny
txhFwdyJK0fiNrXrkPCLzb+1WuFscGBjiV2YSYe9q92Vlb/65qfdhnjz5+V6yjkWBnmEvT1W9fQQ
gMtCIHPTSCdoRpf8wjtyr6W24aEDN3SRQcU67Exge5w6lS114mMfwT9hD6Ahxb7CoNTrdWq7CTDo
N2cAynuO3oLusShEZUUMQGy3AMRbeF2jjWgUnb0YpW4UQ5C6gJvMJGdZIixLvt32KLCWFJ1CAgkP
18aEQPm8Mzx6ggJ6A2WTeKBjnJiIt+ZIhlvPXn3M47KiB42q2Xq8m1M0+M0c9oWgz6lh7apBwIlT
6YG3aHWo6ik4R+vfnTSXfKtNKFiFPqVB1LBEFiBF3m1OVa9zjgP/SU2ZpXnsKGmc3HZChdrupdrT
zFS/X4QJ5kiDOr4C5sK25MjI48mE89MqpmOk3OG3uHUTapN4tPErfhG/ZmbiwpqlZdVOdJkIVb2u
lab20zkFmn6uiHxO+v7M/jUjeQGsdKfPowYmw3rTmw7NdM6RQvCxasaEUr7uUov22b+ziARg7vw8
UqHqBx9suWdazK8q4slCrQz4uJ/HwxTe+ai2DTBE84EufpAIyLN4FWaFkZWJMd1kjfFSPz4Z+O6U
ZJ7l+NBkaCYqwuyrT6tJCU5XumNuHIfyudNXDCPbLZ5zNE43of1Mr6rbiRdXXEtVp6QRlDZHkk+U
2GwluNIVnwuRrckrjSwhDYQncojexx3xXnt2GKTVEg8fgS1ht7avc7QY+PIyxJpM/ETfc3941MZB
o5H3RQjpFdXvH7T8gZOA23E2kAHkdWxGbGVDN5uRCDRpscVDd7kbBfpdBNWzpO59DQ3UU26mfnWq
qTPmo0m4fWH+X0sG2JNAWDK4Ygfvko5iYW8oCWLlZHRxEiTFWJSrn6XtKMn7XCG/yVohNs5Igsun
uoQlGBJWb1+O4ote58slHNCGJiBOF55SIGz/XNB6KL0OhNgcwgCmgQoAF6JWwMKQ5JrpJVxOa2ji
4OXxQ5JqYKZwhr1DtTpKwUa88nMQkD3NgQm8FaIlKJgb5/SBIvztfNFB2nwVz7XvfKaWDOWt3VRD
cmatuGdL7zQZmMjCyxbVaaT/eGqm7SzS6KIHEGEBFH7QrvXw7a53KXpO17EnDXaGHHWdSYlVyL0Z
Pd8SJvAGlGSCfhH1vfeq54bxyTnZFHxB+BJODPgasPMmqBAi4bPO3hG7Ha5gVp4YJEU9i+d9Uq84
SHG47hLbr43/nvRx/20EqYk9HmznKPEPTWtkeHx/ela9rc0WlT7T33EOFIrofI0nMbVM7M0Qj3Uu
zdHvcg4/3LN8Z3FsNi/o1XteG8cfrRYznCFGLrmh2VZ+V1ninV3XV9Syuy/2Vy+gsqPmUmLE8PJW
d93h6HeoRz6FZGX/YGJCfjyVQ35L26rDiQbcPv+bX8eSB2B8bSnysRUSxNsSnPzDays8Ba8paod6
2qws8jd+C2876GwcDsBIKmuLk12gPMZdwWBAZTfLmoo17zAn0gBzTwiD+Q3BP2dbNa1LHHI9W2Og
1g6tDQTy5Sg/Ad9h98/1z28nrECDPmk/EoyhL7AI12wDgfulVYf+b8rQC/RcEUP/05dX6671XFSz
F+j/JwKDPc0IylsE4Oz8ehnASuDpMUb9r3QqF80CIZWNV1F/bP4P/vpteqUyLwl2EC+ZsNf06D9Q
dbpNRc6729NVpgqYOKDcmx1f1EFhAzpmr8On3P6Uew0n85VkBVrLcDRhWsIkzdlmkKX0TRhEgpeT
rQ8I1P31dn8wFl5D6NmmIe+W6sP6TNHdVaEy0wNQ2zmDm9s/OfxQ4N7QNjZJ6jfj2VNsoGsF/9Uh
FZoq12OEdMoYLgVMGKUOoSptneNSJ/6vE418kV+fbwRj4z9ch+UNCEnvezFwTF/OtpYLiOx/H0sq
wurPnUbHBSWEZwgz9fne5XVFHICb/PD5JkiQCivNWW/iDYrqdxGelBoHwZXv2zelF5avgYjTra8f
Q7IVbf0T4O5eUh+4+sJ6gTY08jI/t5Q9qwkysjPfXiyvnIhqdDmwd5A2Hq/TVKdVVdPO/z5MIgTL
ZA7AemhQghE2ZB7Lp4epycHFvW+nUUD2ymg5Ke+hIojt3a0yD3Sp8yMEMMhzl33L6XX6IzRQ7bVX
EiKw6J0EqRtQFOmVdM6Kif8bjZfSvxjuKWPYq80eW2V68RreyqwwycVAhoBQCSxAZTBh5Ol5+JmV
rEA9WAmmdu4E2+YSHDTJvgfAVOWVs8A+h0a19n4aR4IJF4J0rs6qzSH084KKjYTmGlkGw3CldxuF
/qb2+ezqMROuKcBPksRZPTGYGlQ6KeBkqUPOU5OZRfQ8+KTWvOqZi968bdg6CCtMFGLBAQ8ZUJNN
8Yv56Sf0tfE/Ch2wj/Cp1OE6YKtzqBee3Vln+MUfXYHTwNk2xkdaC1/u02Mx3cgWiX5vngWgt6oH
gx2ipkv1b7nnjDCukIRBlVPmTKWg29R0UsUAtAy4Y3XBpRf6pBK3erPTwcTwL9ZQHqbg/XLKegNf
C4ZtETf0lx0ugQjhWGPlHljC1WZPUD0set6Bvkz0vSumj/V5KtUpL06yNTJ+1rGdDTBm5VDj2NEv
c4LV0h5Bd7bht4YLeIlkb3LM22GOM0SdRxyb4QOtiwyT3sAr+ZB1KDNeSZABsqANbhthox58oiMH
TTC2z/ZUVVYC8npsn840nMpbr9YTgU7iOKRNoJQpo2dN5uVmMEd7KCUfNjk3UgFF3WPqeuRi4JtP
PNFYgk9Jv9wBx8wD0l9w94W1whMJdMsGzHlk64lrOh2aIh+SKf0lJidIvoRPMsvNM3vs29BgcX6S
/NIPRzTGWVUoWq1LMpTWz4UYmHWOgORCjCXRerbyQ8mDLKrcc0Ru5XH9BFNqAPjxnH0ZstPVnQCp
CzofHKsWuod56AGoao4OfcbV99tCZ8p/pAxnX+62F27S3ndrydAgM1rSRbAFfxCFNSlmQP/0KTO6
QBxmdBGdIigpSCkXhe27QLnQfS04CMuMCxF+RE5NWmOxNTu9qAOMBSskAWVIse//wMVED0G7P4Sh
4+fVTcmnmr23IUAht1mZvV1rjvEnrNqaINX/nnoNW10Pj9+v5hlYU8Ec7S/pSEnkddei6opCn4H9
dcrJXzvoG/38797yAOWIlUoFHXWu/C7I9woRQf3gGiBwU/sxB2W0ZsiMxxuJvAf5lOJ5CelP8pzV
hHuIQNTHgdG+p0WfMdPvmXy9JqQptkgjupCSzvedFO5q//ElV2L8LDzUHJJZGror0rKCnrEncOJQ
YpFHmsMKz/y64PuMZS8Vwsdfug765yz8A7x5FOSdrK9Qm1VVkTUbPKfSSb9AtIlrydAY+9CMzZT6
gHXF2O2LC91lhzX2Uj6OdVX3s69498fOq/6lCAk9I1WjxcXPCKpWyTiDF9w2YB2217oLXDEljdC2
CiU5Xwdufs8KPiglMIQFatHMkK2m/tJCoVNRc8l92i7o9cvKl5fiKF0rLcl5om2JvO7ASIeb79Ck
f71KJH8zRdc5PbL1Bhu6JG5N1MVm1T9aGpHZ/2ioIUC9t76RINjt/O9lgz6PnPr4NAaEtVPgzU7r
/gJulvgEHJIX4G8dZPfPFteVs8pZ2dCcqO/92uEICREpSGH0YBgI+F8I/040DQGQvnFcYW1bkRjs
XjzDNPbqPvaI70VDpDI7owPtT/7EgfFsymG7iVcjFTCFPLMQmQkbW/IBqn8fq+QsbnFbvRz5m/PI
TcCNFaWpTVds8pDR5Ne1f+WWPdG5FNi3yKyzoYUfa6OC92YlPl582d8+Nd/jSdIQgohad1Jg6Tzz
tFyQJdS3hySvqzppL0DyALNebE0P3PT6wQpnv2lXeorigY+Se4TZpaQ70YrAP6PV5NpbPTYNWXif
SqDrFQjK3cHRx/arRUPiMeLUzQWSQ44JlGPv0eFsbuxtx4iCPjjvUD2Y3cYhLJGWJOMlIFnepJ16
neem59hB9wuMFRjlem3VmlJOYxicpLdPiv+MBeORP85UwDzt2vpZgf5426Diz8Jp1kPakDVTpb/P
QXq+DCnPKaAfyzRhl+rcrM3/4gUzEkZdY0BtuggfHSnpwojNuyZd4IzmgZoYD2wBC/CjIPfau+MF
/8TOjdAyQYIhasdKHUlvnq0lxmQ2nOfxJXJdarQYLqycOqywRf0OJn9RxZ5SLg9ncJZe8WECmQn0
iWDqc5EMT8qIfQYOL+OMaW7Ptf5OcHTuZ0gStbQgcl2l4r4VPYAzVa855lUO4QCSYchloUKfIqPk
7yrEEv1f8SCBf5Wb3G+LI7CqbxPn9SfVBWo9eMnomvxLqQUljxWe6bbbAAQICoqUHKZb0xh2i6lU
okaLfTd4LxecwR2n3vDja1ehjtvm5TLiED0o4mVqTEq45Q8yzibeTX9qyLFsugamH7j2nm/9ZSt4
rDQcVWaiHAmChe2mHppRfFazG/VEuiQK2XKxt4vaSK73VDlZWuRemcuGEZRbhrgDvmbEruSsvBqe
4m5f0CRK2dZHxPLeq8QB20f6P1SA0sydmr3++iXRom4RWSYr04+Q8Hsy4rYpbb/+aUnjpp/3bWDB
zm/rRS0DImbRZp+vbb9ujL31B1GVdBRngqh3GaQaIphSQe2m1GURV2jZCPA5O89wjOuxOvrZ1b/N
j433KfIYelox1+i9rJFigd/CXjL8RUTQd3DnJ4ma3hZyRQDkdIwrtaXHNMIXLL+Opa+lSmYsyDdu
tC5hmPsOyaEwW9fmR15j6VOWWJXQOu+YkMMf9rF/9Twwh1wLwsuyCaFl9m1Wd6vgKgHM94ZRWNe1
4T/aRZJ1Vok6DuUNN0bF0ugL844eTnruFhipXaJYP0g9ccytYAKJZHHPuVD7v7T65LDTpsGP6hdk
4W3hO6pmGTFuBwKoEqPfCiM1dj3DvN/fsR7vAuVABTijMnL4q+hC7rUUYOJ5F+BMK/6OGcH/VLtm
j/boSLzwoLfdKHeHJPOMhLGO39W2AQ8KyhyeW4S4IDrypl76JP4e67cApjL4+p8OM/Wq/y/VdZAw
61gNFGq+f5JHUIoTpxLC3yU9C+Bw7gmoKYrQyVvZ9p7hLwzQ4QKVk0yRIVhOUg841Uo6q5uOpCux
MEWsA8iYnCPijLPnVtctGMBxKGHbRQbHABHzNquJYcLGj/NDvwKF9MwOL9Ls08CnxWXPbxX8pNQ5
WGHcqzVHrsNdsJbUvnmgWHvVP4N/sPDvXRghhJPb6mQgTMwlOonI/ptdiGCH1sEL9vqoQMR2xM6E
V7zkbBqdcaDWef6Qrfy/NteU+H+QcZzScz6nGmRqMaPhbAOLDM+Trdm8Qwey7uc8p5krRIIuUOWT
qAmsJiyelXQcZ7X7NVHuYubbKfFMzW0qWaggpVjMZPlnixVh09A852GxzLDYuHg/Y4SBTYfK7hv7
zyEgGbAVKvNxVYFZEKYneCwf2etHHdBBUqsXH0EbM+Ec5R4uyYFaMaWsmBzGvvyzLIRiqho8Qmbf
coo9J1P6MPovMF3+I5AmCW2XRasJjJHILnujnq4aDhFFMfZlHo5cjbFZS/doKH2vFTMotSXaxwgZ
Hec6MFaZvFpGJ1Y8J4ESoiKHn9GLL0f6j9peWIKuh+bUwepd+BEzE6AwMlVNtYVkMRXqLsI/oAlo
zXEc+9fD3w78KVM3lXqDGDTm2o38ysy4o9ZTN5r9cj6dRec4tGkYsSkOayOAzGF3XC31/lXR9MLi
upzpCDTEiphW2rLJnc1Vw4kKxHwyd4LiRPSHjcujGl19BPRUQkyG3ssPzVgGuIbJBrY3S/SOKh3J
ZXVBLZrwfb3FpiT+To+6tduzEPvdJT958zPvBRlfYXgHrotN2GrmQx6rH/98Kdr7+IyQeJd+Lbmi
NOox4jNx45BTtiE66mTZ3c4L9tMVIb7jzXR6DdQIHdXD98NkW7pQBJ+VczqJSHAjpUa5neM1UAqr
ip+pqFWMLz7Zm9hum4XrAzsfrcUQlsga900AUzg9l27IH63BH+/Ya2XZu01aOFxEDUdhzHyuEqBK
r/sbeSQXnMrkTKMKRPoCytyhlXp7LXmc7R6pstpsPmJ4XuukwNKx05bVRQgDjaJ1TnoSZeSFk+GM
ZSPLfBOgRsgIBjImZqp5hpu9hRHKeZCwYqbB5U1NtqiRfEBYQO4lsD7+1cYeS9/X2xR/5LmYVa8L
Bx+FEpjjMyjJ/xwfVcebwvuF+KKEje5PR9GbhwUwyKEY3IWWT9xO9Y1kCWXip3mo/A+5fc6Gh/Fn
6rlCm8jJ5DS6XAveUyBgTc7j/1K4jbqNeCgWSfW7uPxOFF9yfeGSSeoeskdi2CAbBpTv4VZORNGa
We0l2QBhgzQpeDFIMaACXyqdaixx3ISF4pmbliTH8voj/ZN9CSwqo7sAu2ZMNAw4v4iyqhEbzUrC
+CPLmOcg9zK8dGLbVFfBY/v2YeZtHp4s/cl8Tij6o48xscyOCriaLmO2GxUejoBYxc9n6xqX8PkR
22I0g1cbGOY2iQNtQk6giVL9usoRoHXeaG0FOq4ypdROw3lyu3PJiQsia13oxJifDYdGDxFfR2pB
VAJa2hljWKpMQAJfEgeDVuVCCKu5suB22seCXp37Mbbd2LATunu44QV4lkBDS/G+jqkoudN1XEtX
m/rheVEcirW//DPnqlit35fAtAvOsyKNe8oY1VglUi5pTctbUAC5cd1EntvGWJunxM5Aj/04Ga0d
wAynR7vgfBkU/FlUowlYgtxesuTlJCf/ezvT3CyxSeJwMvMd7/MZyMBG2fAJf2bkK7zCnk0oMFiz
vkRb+AayGPNGwRyFkrbeCgIxhjT8ATK2FxZqS4cB1veJV99XVqF/0sWBIjl3CV0DeQEzP4ki2CdX
19iUtuJ9KXqXd7L5djI2yer49Sm2yYGcO/O+SmY6mI+Corh9ocfA+ZR40Q0MWBY0+u7gRv7VII9n
wp2/djLtWTiKF74+cdH4f114yN1re0UaZX7tLMLGxa//XDBD2NfJuu6wfewzW/2cY166vxryP1ZG
Xq34hkwwjkp/tzLwW+XMynRDALOV/Oq+1/xwyeZVqhaycoRRAsUlp4gR5gkuhFasaicxErEhYo6j
/a3hD1+nVIuigyrv8X1kCn+XTNAnIrP9WvMdOT84TaXit7041cHxqxJ+2cNv7d6M75v4nu3jIXYt
lAepIgpdzjZhU2Lq3SIyD8w+vitxFbEaWhaNnIw1thLdyTpSby8WAB0FOYwMh8TOzcqdx64iCgMT
3CuZAH6/4h9FBwXdcTB/EfECrnCifuFmsEnrliwZe1tL/WKn3nD4srxu9e6NpmAdLTWVjcK0bsYN
khlVaip4CTpSyU6jw9AZ6ZeHWUTHQCWDP7RKJaKQ6fmUxWDyEBnKQHEQv8z9fUy6YMextb/b31eO
1KBdfkOI8eySnlGZy486j+EPVLuWwJfo2A/Cy2ji4YofZJoSe8v6N8SVJ/Yu5SzoyF+4Q7Qt+DMQ
MqLDQsWlJkBPnSKn/uCvwZMfMQUt+vZ0TILNdQwPtzrJ64awznIs23euOoD4Z0J/pDWro3OPOlwN
4i5NB3w//KbXr+H9yQb5mwpLJrOvtuk+cvzwweTQ8gbIGw9tpQAMB3Lc9BWSeCU7+OqOdWTYDnox
73zp+wVx+WxkYAvoeYXjvm6jRLaHVQXcqh4iZMplU75vmgxlQHE1ylbJjGvPqlK4yjN3GRMzlUAI
iWvDOHB8kNdiq6gCpCt3wTcQNUAEdO4ZsVUGzxAKBfAR9NI2jr05ryZqB3M0/tPkVNznVGXVW7aw
VVcUbF/DKbIEL/1XbqZxsOi8z1FBRNJPiavx5WEUPVEPpnYRzBc0XvkPuikRbkIzen73W5fhClNF
RGKE/iMpSANoGgZ8b6XFv0lQk+6znGap6chDxThrpLULbfNpuyWaBk9hbn1U5SxZc7kZuveNF0d9
n1/ChDdF8KxiauTVAfb0NAfLem9ARtVgQaJovHfDXpw6VogIq9zCGgK/oyznyzI3hFicNnxaTUx9
AnUrEgeQMkK3xpmVncl+eFgqULjaOugEnCuPwhc0ANdu0CXzwQu3wjRxwDJWGNccfiJt3RbD7YWx
Gs1B2skblRYMGzIqac9GdJkY/k6hXW+yNDmC4AnWFpeS+cO9oNu2Pm/RfgzpmYfUOJ2Lai8hmKWP
RKH3cxNS2ZLxg/dJwH/NaTBjRQvG0Q0/tqaadtuZFH7VVdrO9yc0qk4FiE2afm6zjdCRq17mCIFH
TOvlRg+Dbw7ZbF+RhSOVNK901KaJbso2KXeOyllkJTfBi9JYND52b8Aiffk2m9e5vuMHBoumFO44
G7zNGK9qIpQSVd7YRSi2ycMSVoGR7a+FfhpkOZnQ8eb2+2HMCeI1dgNRLz51PYIZSmLv2Ijy/af4
xNbLiMmGsy/+4OtHYxKAnjbbkZge5fHqVKnCmlK6xvL1ZXX5bQwHrOeLyv9aJbAYbzCIl5jR3fJu
h8zk4chCN2j1FcnJCxOaN5mpFIfZNTbr1f1D54jBu+7egej/jlbWIRFpMDTMY7z0D3yaAyC3tkTK
CRlKUhsyNXHCYuCeRzGgWYpo0TvRh3u9kWS1iBdntPTKnOeovkU9D2gQzZw0nkKp3CjdQg0v0QYw
B/Um0IeWT4MftcUwOaJi2BXYYD3PnXoK6m2YLcKCO8TK7lG+r7ZomD+1X4+ZxAWSwu9GRYF5tHQY
Takd359doHBnABxUAxtap9ntGx8m5S5GnTMglDvTQPTgjFdnWXOGDF1cbGrsgvN+LjRbM/bJ8FfP
sl0BwnHvS8/15p6CfPdP9gRmkYrFVFlaWdtjnpIn8Edemn3XclLC8Ua/l9uMqK6Tit4PF0szsoru
xClS61PFLfIeSFdE73Wh6+XeiVsCClYKpBsYPiTjmIuedcyLhXPXtVcUVqJ4nuqwdayW0G/FCMRd
DnRZ4DHPdlaa/psmGz1+8ZxLptj4fQokFD8XycA8g1eqW0iGvbXlXm9rVAl5WFcdSwh/qlLlNC/w
BYFo3nFKSIFKcBoeMI1DtpAyN9bKENzD0M576OgDt4VudF/rPc9EUrGqs9KKSDpsxCOkw7Cd30Ai
gR8c0E5vjQlXXDQkkBw6MIlDie8zLiOsJT2oHQGHY25sddugRKjqh3SRwDlxwh+iYi8DZ5Zhe9Kq
Z+gNFGDfOSGvEbA1cBzo28+OAU7fE7RFO0LNEMz8VUuzdqg0yFwH//+YHPASrErV1UuvElh/3iW8
kgcNpdSITV1W8jzGo1Xo12mmDQj9CUi4f+0r+LOMHVK3SOhbsJasrlI8PJqFJJZaWpAH7X64BMjF
++BDTaSfGicamOdlOYKsDDAQdymxiQ9BLD9WpMiznFThE3+WsmkX19R4e27lpjbp32HKbAUM9stj
8Bk4F87b7v+8ECscr1yh2PmnCLMySfxIwcZH2nBjUE0w0YbruOKcEkvMjXNwIuCIof4gN4ESFgRT
WVbSEAWvYwRxSC7YkN+2+Kc8/eVsNc7ajBeyRNzbeGYHTReH+7rtx1iLFfJMTc7EMNI3qJbVdsOC
kly3YoEYh/baNJ/UfaG+iqY77kCfNw5xT8Nir0nSRZCYBv3U+l8pCKRsbvwS0f8h86Yu7iJc0sXB
v29U65gOrVqgHRt7+VIiNIVNSph5COVkf906UALWniWHZtCqnBLok8/h9OXrxtLXWR6dCRIHbX6y
SOtzbAYkPxNp8ejF6Kn4np8dqderq89Dci0VDO2NtldaO9hjLfkIdpNjj4r6zsi4h9BZxRoT6+Cb
xlKARZUHswOQAG0qu2AppXl98H3UQajYz4m49VAxI/7K5WCNY4r/98K8LjNwkC4hzpSHRsQduq+W
1blYQRFjd0Lozql3w4JW6rK9eOtQq1X3uOI5/owUusGG4x/wF9rYYuDVxTwPEDvlzMRAHFwYyZN6
fKB5bXMY8dJzRXtG9lHKCoKcLWruB2ZitIVihFvY6MPEjhC/rki2raI2gHauzGQN3i0RQG7vwjWY
JJhgbpg1mRyqz7zvP1covciDbZkf+C0b+NGNQQXwKW9lPavngQLgeNdW3jSf/x2KhxUEh+xm0xVl
wyyOhsOC1gyJ1l3EDB/wMGIFrwAQm5HeGUcdXr09eqb0d1XDW2PaKhEoGv0JsNT6NadKJVGi7fIv
4sv9M17c3x5VzoyeSvewBn4jT5wkeEP9BcjjBke8fq2EHfs+uYNhLnwQDrnIN4vQSSc8yLtOYAxM
QzWpYVD6U8AGsWKUbNgR4eJu6GSiQFeZHkA7aH4XHpPglx3CuE4YaD5q08Z/g8i6MJKS//8S7jE3
znmhVLRea+Ins7ChbIZg2LKHSNYZ7th29UzOm1Yc8mXOb30cnJ1xRdqGE1rIg57mBHkzCU76lJPk
XCYb1gKJedcGOmYxGtbhRALamj/QgO5RDFjK/YYuNMdXhj2DXrbPrZ0PKI44lnmE81qDkVshLH+u
XC2F/EQQku5czz/Vz+Fsh+GfjrHcjkLHQliCqCqS9G1I+Mp7KO5K/XoKvvknnqbGhFy915licg2P
sbsywc0iRlrPOu9docHGniR3nzjef8M/UwiLpU3+AgHfBFuMvVbP58IOayXeZumzKTPMNaN0GbES
VSRiyXUfSpMd6vg7lSdz2Jiil9dQAmPWGEoI0eJBR29ydXOVCTJPoELbo2eKz93xLi0QrIvxG34K
iJ5FuR5EueoHvZxborOFZLI/BfmtYMRTXWkpgQhYOKtfcyCjALeHfoqdffmcEgud3b/Z87FBWUq6
h/eidMAjTqSr5C0u5OM2Aje2yT87UXaIBVb0r5PAIp0mGV9zzhpjQaVp/eQY17AQ3rEYGBMOh4H8
k+3iTE0ssP470qusrRVbag+LZClmTfHUD5Z928xoH4k8yuWKHZHpgHxhEl1xCauBhz94LI6CotDA
B0BjjKzMJzN5o1px6ykrKvU+5J8ESuLubeB9+b8mO4Orgqwwo4M0yxo01P0x0YSaNcq+u0cYmBVn
XC3fIwO+KXVU4dIlwml3cQE9esZo6zJCt/Xgro+dmyU9wFerO9R1aleIognlcD2dTvsRKEVWxKE4
CkqCDNz3CdQplTharVPREUT3nkZv9UNGGCYXV4GjtfACkFz9yiy76rG780KPLI8Cw8jUDwwL94ks
1Nt3avqRKYb97sz3XD+vQ0rufowva0GpTuShOhpr0Z3InZQIqCn36K/SPqcnzL9Aw59H9YLdMoAY
zm/tEQnBnWMFLp+ELN4ST7XKI5pYAKDZFyNKV63mXy1lpmbDhFSww9SV1v+uRWcVnfqoPXEv4WvS
vhXjb0M5rTdDLQt5j4zjkYMKFNfJD042A4hBlxUutDh4G0R4BLzB362SkI9v1L26NQa/QdMh9KM/
UbVOaz0i+nev2pNeXsDmDmXGRTj1nue/x8x9msNQZMsxqzewAT20LcY5TKAM8h8YjbXxA5FxJSwV
BWEukGQ4WmsCn1sHK0NfdNQ2Kel3vY75UTE81webJvQfzLPqw4zy/EVKULmuh5S/joDHVxRfFWmZ
Qor3r5Q5iDNT5iuqsIqeziRN6h3KWOf05PvPpP9aCM5dNDAagXhxu8DyAoQm42ivVbBhOsZMcYVj
9cPE4H7y38tm+phAH9p6xMZyjSPgBProeutMWGFAubuofub0zycry2CiRp7Aw51apwwfgjRNZmK0
7GzCrjaq6io81H1+9JSN0TuQ6y651R9QwFgHAuTzICkonMG/qLI5BxLdhkMMkQcNn9iEBnhc7QdF
Ntg1yDulaOMpM1qrqk2y8mNIv3WgrjfEZQmun5S4lT7X1yjktvtPH6nGMVYyNRwVyrgPUOz7UqXz
89DMEvu4QZ1f8e35mPoui6o9st/m5QutXCPPGRfBxz466C4apkpTMGq1AIBvNGx5rdPrZ9BrUilU
sxC6NUv9W0GAv2s+YJ7kJVKvGECl1eNnMlzbz2CWz3CfoaqomERiyJemtHrTewbLxpnU5MjNreb3
KyhHARsJYPJDi9X9qocjY2Pzt2qhhsMd3ghksIKVxY5/pwFvWonK3smG4uedzr4R8t3twPn5pN+a
/CZyVABULDaQv6SiXidh9PTSd/1kp6+r2rlW2xvzTb0VeF0/c0QRhue4dTVioDh5watHuQ1bT9AN
2tLsrkyEJYeaJc8FZBneK6kGqUbjR4nkzoLX116U+GZ6Su/5EnoAG++5lS5RFSA9iU4eZ1b+Eg5k
JtakVgAzSg5c1JNLdEQdMSw8ffUhNkBduVRTxlLCisw2OzSxuX5JvEVv5Tq+tIoMr462g11WZfJh
LGPIyyeDP7ufOU83wh3D44lL+gJD8bChKq25rzgq9V8EkZhTCYiu5wArNDgJRUEY8r5QiMnKU7nP
a9yuPAdqB0GX7SmN/dQdKvCV359wQRpHI/6R7xwth950HlFZJ/aPbsCoLoT6+yDhZxVqpz+zXw0D
JV4Axs3s0WPzbLKIyYV829Lhr//vl3q6GasXoeQmiiGu7ErojvnOGfJMLj4t/9ZZ3JorIZIDcjXz
Zug9spaOxm15XNHo5XYWz4Z/e/pQ5iCTY7O7BcI5Ll3+q8DH0z25KjaXF18SKqNKsRFQ9FmSLI8m
lFV2HWaDi0PTHjUvMxl8SRkLS5bGfoEu/cB5kxqaaHzeQkxtZ84ViW9vBNLC54ku2sZhPgw2AcBk
ScvLDF5QEKIQ5c1ANHMGW5a5aQ5qEipzScL0LpegMY45KSNw8EN4fU/D4qpXUrPREPgM0yfj5NzL
buPcjH4tK9nbaGBMWBo8iEzRHQVJ2HFMHPUNbVakvh2uzXsO93tRv8/L7DjQFJOHYFIz7UTx/s8Z
7JbBCAoLfirOcqzaYlolsTZonmYPCYL+9MVw8BUv1gqeFVb6UL94dsmAgD3gVlSzFo5ObHyIdVhI
RFL4u0/PsHmgDAAd4Q0xZUNqXF6rU5nT0xDoo/ujVrjB9K6CDd1zWOc+8e59SoZerTiHMlGrRXHu
52FU9a3Gno0ozGFipuGs44aJDZ7VvlaqpV1khz31e4uGjomiQKHBpM5juCL0KaDE/LhuHQ5HpOdk
4EmA7drRIF2GT11b0iYeZBJq9sfeIaRi1jFkZBL3i1QTGw86NMGr0XDEqyXPhRRRSPEuCCrBH52Y
TUCRcxNXcwoiaALiAJEaGFHCycSyJtFWhotZbDT91HUXbj87m8CkQjpD0T4LqbJS/5xxXgr5uJDe
4mNATEeqvJpQpoeODxBTffJh/xfW17ngPt8CEWBrrlPx2cCxLN9/3BQljJwkjc2kdgooJgr1JQPN
p+VtFgB5ETEUKNTdsthSlLyL9guQoDPokdUqdNmgqMepkjLIIleq4ywvAxOB1ZNp3BdxuQl2hVv1
KGa3f8n2K7uVH25jmkciFUAfnrxJ23Wg9pkL7Xa3WBBLB7slk3z12ZlmGUkstbY/WPY5eFAg/+LK
XpDPYuJky7unTZHeEbceMUzlj734fybEhWHRVTMQ4hEKDee72Rs5encb/0IyitpEl3BHxuBa/ZNH
17ZIa3NUWmI/SBALvbOSy9d7iOaDzymJW4+6I/GNEtTVQ4pBzhoKENijq5v1L8KoZZvrg9pe8xzk
lKnJCTujZDVJ3mgh55Mex+nOj8u9J5k5IcWisqgqIV0LtG5TLJbV5szCQMVn1Hn6ipCeQ1Xojos5
yiMy1tOVz+DWxcfAqzjEnlmK69ME6ErkRMMT1t3JUmxXd6MdZp9w6l2Ni2RdCiPwFXTTa8J+vqHm
PYmGcS1UH5S4CwdDYFRYiv1Fl0ZSub9YNnOFwkW80njkZNlDZfAVnLb+oZkstmdUNu/kqL5+N5+6
kZ9yQhTdMNQHzcNzLsi+WrvwSquoJBk63D7bSyhs1zOd3DQ+Fhy8AabO2s+6lOzAgMT7M2haY2vt
P8x/XQbirvoYCoNX/oLX3zLzzICwJzRAKT2VBWt2ypLAc88kEpjCrPWojUPFatqiKJT/OAaqiFkH
LbjNPI+0KwMEHH39lREzZC9eGOzs68iNKtHWzhlDzYKwz5TAoAhRc8eq1C/wtmF0/wufDJMPyQl9
/Y1Y1mJGz6n/Rf8RsMEj9rshcqlIgkCikVSo57QAIiDw2FLdTz3fCRo7OTbj5qRvpITAwIs3Li2R
nXZFX7qbySZOn0aNGckn+oMwUlhnOle+vLu3qrSFVRumttv8g0GAZG/7Hge9Fi2k/J6OPewK0mdb
pxwCmEHh+5F2HX5Pml51hH6w95iVCs6xU4htCH3mRcwiH+VzBdhqsmxUAC7O4LNsvkPP+TTsKnd1
TUcJwMA4Y6iBFaG7ozHb9jrHJI1zg9u9DcYDgAhTeHI4/SWt2XQTpDD1qumRVwUtNemV2eWyHTXu
aLkQ4azg2aKEsJ1fryRkWUAcsQIYna12gKRk7+hsc0olFI9LyPGlKi2b65UX4eZg97gfcuQNBppI
IzN8boi5N9us4+4qCgn0VvZ5GmGPBG27R+WNZ3xl5kRsq2639JziZNTQJR1NOkWLyby9xdqf2EeE
gzfiXSNyYQ1gwT3PjWXV31QVBmpIaCyjW+ip/GXtNiWAjkbw83vCS9ck5k1FV6rEGER1TZWN6ng6
5ABs6b3gGljZ2QlDkfC0cSDFHKbIOkYdNszWEm7xcPmDnjBbPvCOQ5iCUqKx7ulNyDIX9y9Tu5V+
ThH0b8HZD4ve9Ne3Cq2TlexVpmNOvaPscnon7LwuPZNUVgbojG37MXaeKxZwDBfQpI0pS4X5dhoL
ggNtOypNNReOYH30uDwwFF/p5BuollHYpGNM0/RRkvsiDI8fCBJYi6AQEoBvxdczED1A5oVyBeVS
2MxH75mf5SMJHASRGqakQH0dZb18i3WRfTUwq0eliIsCqpTTlGtaVndNjwRxQH9otzBExNtqrrIS
9UL7iV02z1fb1hDWL9Glj9mftQWfLH+qkQfQj3QCJC2UoI8dIveVfXc5AP8E0zSl2Eo+DbB2spSu
nOhaUekOx8xmFdEDa9mmihl91vT3ES7hozncal8AoDE7WRTpF+nCCzVGoSarXptYj777tlTHRt+i
SMvdG6fw81wYVciRWiBN3l8qHeJKPqgRCzO1i3l+fd93mAD/ovqmTPAbXuMnkQsQMZ6fh7CW5AA1
qwDAgvCpnD9OoLKs3VxQIycTdid98XQN99PDlN61r4UBk7CLcfil4qwU8fvkPz9o6lUFp01zUzFn
jjPbiP1AmwJTlMbreXX6aYVgGrVgKBqFJ2NX/oToNEAPG6yCXFqvoIzBqMhyZ9rDzYNIMQpZ7heJ
M/kQXaEQdo/gVKl3/93I5KDCkJMH4e43VP5/P1nlBC+ErSPtcf9sHTzF+Nc6aUoz6z36sBbf3qUc
KRFj/3BLEfOzfb4HoQf6+szydzcm8HnZLbVUqy2cw7C3cLJ1KBfxwIg8R6oxzd39bns/ri0YBwGA
clrNpS6RapjgNoYvQvvrCcBX/k6GRCpR+e0N58+Ki099SJ43G+JDyEA2+KD5nRipPxPPTSVGtQPe
FICa7zcLyz5PB4ACZ+JRKVvn80NPWOBI43rEViycd3wHNIfZRz1fKYDrYtqx6VvvFGfMlFpLDa25
PGPqJqtR1M2gRqMJIyXFJ4gmhRWUx1YDTK9MYwZH+EQdogofJIPTZiN3ATExi9mxq3hwa8A0sxwJ
idFNDJdVB6BrZ8XnLeREc7jk1JdptCOJLZwUlPqPKZcdssMf0yulHMAWqrS0Q7ZEj30+Ditun0pb
C6re9u5j6O7/dNuK8KItKAzuwJgXnXD4hkFnyaQI61CRxr5W5My24RDCqlr0daQN/q/U9hmgqm2C
ZJ9hDbl55MHYlz99LzMxzhidV9ymYOUfe1XonZ+h9kmw4IxeF3f/idnR1V0vol7y3jrjKGh7OhAW
rjSkjvSnx/CdD+T6T/FhW+Q+arnLSZqfeSZFgwQvJwCv6HRbf3UtCbrBNwofrTvFh2VrDgQdxfY+
Oa9iAP9o9C2LRZ1581uOlE6e6pNaXeY95hf5C0ZRHuI2jYcpoZ3FoPG6CriBrr229msQM0hkRJS+
y9Ptq6tjX7GWO+Gbhj8MO6c07wCbpsr5jLaljE5nVfd5t9vXYFUxalBtiXUK6p2E9xn4cJ7KNeL9
tBs3QR9bmcRRkKRvh27/gtnBvjQT1LnZvYanA+sk93cfu/RrdaAVDoukfkCAoygyq7PHCbYNdxLC
vhJLBrNvobgqDTET1Jtc2w2f4M7IIiQVUU7BEjmXWN2fBWcqSHQrtkZU/cCsHjtaCr/xvD6XZb6Q
FeEx9swRiQDLbk7wDLaphBTDvPwWk7T7eq9I9mVdZMT4yAOmX9w/5S+NUw1OWoa5NH8ncV/8wXO6
h1rtSE3y/4ukgsj0XX1xyzC+dUrJmZ/e24Pr8dC/5hkgWeDpqW0WvBYbEg1IPC0/HRII6/TDazqq
/5VfbiKx6+RvSA2NcpHSIsqa+C+Kk4nR7OcIpFScFUEUqL6+MTYylbqbYNupPj1ka1aYvOVGAm/D
wYDTQ5/BFBENw4BHLbnmjGuIk4K0H0aJEAasabLajPvN4/6pL1F0Xte5chVlH9Zjj6M9gDArzezS
3HMj7yvcMrXg7UihR6W3rah9Dl7tnTE1hyoE9TrUSIgExNmwcolTvl8K9EF+w1eCjlSi424YKUf9
oEjmKYLUBDQ847IAPdrk7Iwcpvh5DpcEuzagaqtMjjq3pYLLGGEtQfz8uPLD6hT4cxyY0YKpGUIj
TlAdnZqmZ2SDMiQdt9VRHv53i4lYghPmCnD+gjz+XhEENBqcp46md11v+tv0LNUydZXG4Ps24DrY
N7z8NhdZja1GZNPTzPxca8mcAbztifuAplU951zSHsawp+gZ708pzeBq3oNQrno+CyrQTrQY0TPQ
dQEwiDktkWI2NwSHlNSWWr+eD+bqtE6XvbGnt74XkiK6Ay73tJTSV6ufQ8gO3tYMo6JLRRloMGz8
2n+V2oIK334Gg0Kxy1dpISZw60OIN3oszLilcXHygGOY0YNn92T9CFIL/37kASRpAigDHdZk/yP4
1BlAEH7avsGVPczNJDT4p+WoGTuS1EWo2obfL4/N1Tg89cSRUsa9A3lfHlQQ06Jmbw3wEdhr8KDB
IyyWbMP7zAXdbMUbEPBz/M1NZRTKMv9CslDGZJMiqZlJg51WLckqSIqDlndxhbiD7d70QDVDGSdp
zkgofLTfZ48ga8YFmX5ZBLuYaHmyJkn7wMCe66p4/Un87UuU8caI75YeKBG6sBGI/io/4v6UOUq/
hL5TfxyDOoQgzU75n/znfjcstFwp0Hbb/R+AG7KsGfCra5nkjb/aATwYKU3CXKi+2LnEanoD1KHi
Kml1dY6mNwCEzvKGw+gGcv4RIJeDvcFliR1fyAm7s6fYrk00qSIWD5VFCSlL1kxYr9qSv+b7HnFi
Mfeg8ALQIPWlTyBlTW3zR0Xccu0WLWZ2D9N3petlVApaEFJlgdNMlphGtPF+UY+dGzyZ+Go32s+U
LUxnoPgK/4QEM+vvI+v+rM+UQQdbkDkF5R5lHYjvSl96rc0An7tC7c1P2u8h/vbYHNHQK6+HOQb5
30+gxKOsfFewwt9jTyJUqjuB8CmezpP6yu+Tq8nVekMwDiWljib28CJPcSsPVfWa0KNsyCSeS0O0
iuU9ENqxWlnLWhr2X1W4D1yQlGRqyq6drOWWksuN3bWGWEJO9eqRftLPfu+Ofh2Rv4AdNUcULX98
leyXmnSqy/BLMQMuzwis8ZV4ohoRIRRc0IUjocLAMCbNNfdGUxbauPlSXe+ZE9u4mUHm0DorLrZ5
bwuwSrx9p2ultRmvFzkJlhPiiTICtk0rkN1nDxH0zGzo62xkLH0UMkJBuoCC3vYQGD8iKDzmgmjf
xAafqlXt/2yHToZvOHAsxyFLWQX7LPbA6L7Ld869mG+M/A9plv9GJqIhwbwsOUb5+XTpFlB9Wkdm
dErTNyWoSoFpkQForzaRjya5z1mQw0PNrrKdKcC/ppIFeoVgrzRV2pQCDkBp/J64CpVDywYGmoqr
8RHDWwLWRPQE8/7BHeSw31QaAypvzrpAtHgBaJ4cDNJ2s3G1gkc0Ry1nCXFsGlCerTk3fWNM+enU
Yv1HRDfRsjzLE9v+BkvpdhQKhzBjb5o9/hndjM7rHf8/ivELsCCV9dsLFeAGWjBJMBQ8flyXbsZf
1ZvLF7ZUrSqKYdHJOO68C826da1gl1xXT6zrhLLgGRzRCzx4S0zGoq6OxkPhqFkkGNzDUVhQyrOR
FH3gwnVUsaHsfwpuvGpNLzk+3mUqU1N+EqY+MXm0pfdBKv1qKTFKxH8WcROaDn/knKGIhm9Q5Yih
b9yrqqhCPfkL38HzfI32Muom9YzFi/MGuvgYCRSGgPme98cKdJ8AE28p/cV9rrJT5lvAFJ66rGiL
Je0yNJ1+Z8FcN+V3RnoowBm17HAWoxs2BJLOG87+Vbd7fmfTOWP7cbVEXHBNI9JlJ7JYml72Sz2r
pXMmhbfUGKAfJi0vHsaFn1bE+PGzzv+Mv2YgHAbZh0tNapaA/8pMhgCck2/isoZ25KyGphXBFX0U
3vme9/66Ax4GCcJLjtt9VxjvVT159VfLbRFkzUXEUOewB4x2hiNgv1TFAZJYAI6ZB7JHOYOZ995c
pqmQFBpFP0emCTWSfzipHOH9jbEXIl9Mrk7Te9aTePTOUJRj/eov4GrXzjHQEvga2TLzDONfk6bx
aBZTQrPVU7a6lO396xL+zd3CUJmKlIYvyyEBFx2NAqJnMOsTwBtOmCl9uhsVM9RR9OLY7iyZ8j/5
kChaa4ueQBgx6QmNPT8F34y1K886pTU1CMXmnH/1Ra+KuMVS1hRsyMHOvxe+RkWyVDLsNYqpn0kf
ElWJqV189DIrIGfTnELBk/R+yLFxbD7qG7hp3Mvo5aPHQzkZ4OcpTt7Lu9xVanZ7ljgx2mncLnxA
F2nW1PZ/0ATXn84M1QoWZi+51TD5zm0ZRtYy0ZzzJU/U6d4gqSgITwpTGvKwqzo6j07fJ8aMRnzy
lxxt8IlKHq9aV1low9AaT78stYTo4M/1I8UjhGB+sKEpyyMI2Eoul4YDwOQlnaHbzLIGHURK2YnP
Wp1E4uDHCmhYS5R3sk2gZ9Enx1UnoFFhfuph05f1Sxkl0x3QZBBKpOy0vuAgnXyCJ/0GVqpaNRu3
6fbVNJNr6wQlqoMjMZlTEl5/EhqelIvocCB/HPdl7mfofiXX0c01/96+jHUPCspWts+y4EvJsDLF
zHEmrwwBtNa9PBlTXt0tOn3rJni6jH4r/2LMjxY5ABCyYEzf4M5XV5XvwoGnkA26HTjFU3WMQPKK
6isrvfSAnhhk9vAsbXU/M9YcpbDyI0UIceaOmnG7ThW9B6qv7C1CCHmgAXbTRe5NEpWSstdNeJVo
ZPHyQH6vUVOs/cj83LSy/1xRQz9V8WU+HMF49TpfK8WLkdfX9EaAk6tD1XKdeGxJiYl6toDCd+mR
GjPAgPyjNXY6yQOR1Xi12TvOTFIxmBVmyLqSFjpHEQkh4SCUG0n29IYYJCcl6txu8qoBESEDanKY
H0vmx1DrTHECDJZdNw3i45yAUSJwa7Mzkr6Gp4Sv6yM4g9Vwqk2RRfGsjosa8YLTtQmPHe5mzkP7
AdKkRVvbvY3ZKajV0d+H0fMqRWToIpUv+Z0PIGLndZUltJTYgI+UPNNKpj6wfU3nYxA/GeYsO9pc
QZCFpI/gmm5rX/5btkrxB3U63lPzwHhPKXdJdnpXTSrrXPv7JguGA3aGD2wd+5c7mNjU7eXiQCWa
mE0zhc59aPS3X4+9NlknOyc0WtbML6KtqbaFJnIhkcxTy+ZDQj2kBtMDwTVyPBmBbDPhd/UybRq3
E5MKEZnasjl5R/mKK8dzC3It0Py8nPIVlt5tnxQ3NrRloMODW60ZzHNUl9to/ZvaWFxZvrpLyBl/
LZjFAnFBcCjJIItjqVZhEHqnVMaHXJWUzdmZNIioGEgLBkEOBLE0dlwuYTvlUukq7PbUDXgOYShj
NF2bLP8EgxfIgjtb3KPUkpqeA7NOBvHPZl4iHitncdQyqLjRGxCRlT4m1E/+IX39oJiul19D/dXa
kGHCvDLLFMpaZY1ymg+XlBBg2czkM9lBnUYkwyMWA7WF/bUSEX2HsJAwseoQgrih9w5s+QGvy7ny
pzXJ52gO0KMgB42I4C8TLkm5kDFgco00wYbLyos6md3MH9zEkpD+rZ8PR4cwFVVgMG5uogVheVr7
ly9sLO5Fci2VWw55qVIRqzIKswwcH1qrMy0LzXeiJitu3Ah+DeAzfEvG7ylQ8GDudq8ZrR8ov8mB
S5Mr1CeaZgk8vdQICbnMQnLUCglJ+Bpkne7Qgvm759mF7exfriEpHdkg7A4qFXxrPp0SMhUwpJCW
1HsEInKNlcrS3gh7LgRg2hTD4BT4TwX7MX4Cig2KjbGfcnsBUytzo/bQYvWksL2gkUNWREOVQbzk
LQjyolKu++Q8XS+ix1w5o11sAPzQJ/OkKJopmbYcwZJMt1YE2iwdk0IxDLBnY0Alcet+PfHfbKXq
VRPsQDz9RD6L9CaHe7nPhC4HP2BfG8aJXEyjw1f4G0ecUx9bQFS2/LULcRIbC4E2PafFnACua2HP
MTcVTWsN3Vx8iOt61JX+BRw4wZJshNe8TF0XfYle1l5E0iwXEC51dxoY30vxjrWQlIeyyhTrjb0I
QiRm5h2mV0J8TFtuV5u9Kgz5LqDqwPxPk6vBBtt4G5060whNedkb21u47sDkIhIGV4jorQsQufJ3
j/k0PVxEkE/7scdyTwWRH5benqFIx9Az5VmIqGinjnl/5TKScg/S7wt6nMVCboCawiAW2EPwWuSd
3L0l1moyLt77RmArVN1IH9YXRbK/7zZdgGHcXgP5QVez1H8olJKRpJ9pmsCEdL9Y0cf9vm62fIc0
uGqI1yxGcTIz86dE529gP03D58YjXZgSULuFIYl/2YHY9L7H2Bd315WK4EvvH4rcO8r7YWCIZ7/w
NQT5zs0JdiIrOLJbHdmCYdL+J/icJLSbJsnROmYjOlAXL19cWy4ZS7Wp8r8YgkBj1sFwvavT17h0
fyUZrDj4kxhSkzLeNA9AvOlvOAKVxNjm37cePh6IHrj/5q3CwnL7xC5zIqp0ATeH4EjlxE5vTS9H
ngAP9Qohhih+OLVKNu92SjXBGvv/eNzaBooLfeCNl99C3NbwlqNAfqSaFU8rHhK6lhl5PLTWIGEt
TkFxrwUuUYE2v4mdVP1P/ahgql+epNGZkQPrz6LZ+EgCpwDe8Y3dLyhbRkCq0Rh9UdKDNFvHpi+8
C5UWIo5Xhp4oR05xGgV2RE6Ge8SCUadN9LIc80Udm7lhUSi+AqJhrBND91Kl5JHe5aIjQ+2uahfL
0u6Zj9kFUq6vQ5orI4bpqKuUW79iBl7FUsnE3eK4egR28Ps6/yZurBFDteQxWCOcdfhy47O/ezP9
4rXrO0odMtSrP/G1S5yRys58fPDh0bCSJfFRLs5Q+AjZco6VFzy+BaaG8skekCXnnoPih4NaamvV
EBa/QELOIVpceLT2SyzPVGOyG8cBsuG0491tNNf2RI90TvUXpFHN7Z0zRiOHNJUCz9btQ1E3XA8k
xsfYyxMkQKKyjdSzCAqAyaGNw9hXDfm5oScSK7BTt88YSGejLICGIB7cnsJUpqTFzNQ8N7ZUSSas
2HaAPEJQGfEEra9W74mlIJh+LBd19FO9KLLRUH4Gk+6STyHDC3eEXQryx2VSbpSa1WmPhscxvIZU
3ZD7DgPC+NJkW32AWx0rba6BYDakwKsqsqW25hFv5O/JZVtasSuVVlJphoc5rDtIGWRIskMHkYyj
gYON6CmFgN/jngISsBLVKqHlSnLH1ru7DHnW1e10AGMLPy8Ya509rlyQhkjptLgEKdqqs0noPAQR
Wvmy2NNoqzTvkju3pFY3DpTWtA3NQg/SqHCXBGmGcmJatM72XiE2IpVyLPnTCKosm9nwljDTOW+Y
wZSu06gIM8tGsJuN9Ywuij3GN851BlBMpHujcKIho36IqAq5V0PQbaqD3CqB9im1qkZ6v1BEh5cw
IhEmYIKN0fTx2SbN+hb1IkrLwF1l4ou0F7H/coH7bEiDh9ynk/tBHgrk5Ch3Y9+J4UBp3SGLkZsu
TQULOuwfpo7R2SB3ZrBtR67Ts7rp76Ov2xE91dFQ+8kMjU4uco058lIXRpeEJClAU2stCAJz0VMu
HipWVWKq0WrNVjkUeKn5ynl7kGdDQdvN3C+Ob0T3I70MrEVwFNjFFd2jdzTYbNsY/zZ63+TJSQLd
rWD0lPwO1QWDUdZQJ32VD7v/LVytkuTjPaftNcgpy1TbAtGyJHh04kMSh9o2dQNKkrDk/up90oOq
kS0I7HZQkxYAojmor9tg50D1a+cldujKyERIFRnrPrlFFchRiFvsYKwOrez//ivJ+1TUbnIOL66H
+6tBsgN1pe0j63OLV/Ir0QnUd3T4eQkPh4nNTNYLeBGzbAB8Xg0mhPMyAzBuvcZBOp2KzTi0PEp7
nkxKEREC+cOx1Hh6Q6p2DucVYoBWknFHcDvfVEW/SVxgKwVwP8Sb/b0rf0BnGgAJj4sq+MEWzOfT
o8KyTuFKFgY2Ogz4Hl+Ic0Vk9zBNYzcu8fpvzlnfu7QalvfrKX/EaQr/P4/tDMNQQo90Bcivi5qJ
ZoC8inssVxT93p4l21FZRcYEWEvGjnmZpyZTIrsAWtQEPbCi3PZJ0AiVGdiGEIYyhL/F4GsFgKfw
FYD7tCdE/PJwS8wSCU4naHZBQEwfpGPH1hYxkrjZ86G+69/vTedeoW4fY7tOqNIwsZ0AqLDN8CLD
VlBPLR5Ts7RjtO6Rlrv20itnTlGw8dC8pdHJXu5WMxkVVZnXpDA9imiHSYAoQHg/iL9IQm+2GskD
IVD8iXvWHuzcrWBsXMYEZMc8d/omRf3jSh5+hAopdC3ccwmA1R+a5HwYikrHTqhk4t5k7BGaSByP
Bt0dK4NZIwE+5yDskAoAmS1e8QtMhE8AmcoqR6/KpK2DxWKIHKFXo27FtyGJ/b3xj4rlgeZdw1nO
Y+NakedwRQ0oTS/mv8eRYh0fCUTw52RNXQkiNINPQdKBlXhfaaab75aVe7VTXCFmhHrH6dnRhVC2
tNv4xznUHwz7sPhPLgl9M75c3rtrK3vqhx6MpsRj0gUGhfjeVaGI/tOZuNcttkqnsgrWq1SWPWVp
0q45+Mnko3CmFI8unihity01Q5s6hcPlJQZqlQHIXS5XTpJ7QXLe2TCD+hsmsQpThL9eki+KK4KD
jELeZj39xyMs0GpF4l/wWqGkLC/qPU4SFsqpUizTFnh3QPcJkk2F9OfOwWpKrOmymgl3Fy+Btu01
FPnahQeCiPxwFepdJ4TCkUtJC3xm9xdyoRfZMScme6t9H/t2qicEAWCPXsosw4yRMmFliWBrfsVK
7LpHSfgEozBSyTcp5JjPCGtn0QoOtzKQUOQ+lUmvuXfgW2RhqejeAjjyJ9n7xKhmkr839G41KsfT
+101X4FlXERxS5U5vYeMf1/dfCo0SKpKKXIySxTwWb4Yp+sWKhF7AQrUMEiQBPbTwtoo98OJdH5s
UCjlbJdGb/zJYEY1QvIOia1Cg0h9IL7EALDn4sCe/mmCYvpRDlOnbLxySfvttHsE+NPX0EtNW+T/
I591k3YPh73ihNGLwQNutgIadL+ZLj4Emm4+9r0HrYciOUq4i9GQPwLNLSFrCa0LSgMsfBgSwTm+
HoU71Bn7hECD8yHc85Tt4ZvojQPtn1vGidlpIHNS50gLdoV6Tn60KOx2vxoUXzaQNVjoKzSCZbKe
xOO8qHlsscutoqZfxQm5FqNE/iHLhUTQE13Wtf/0NF+sMjQ74cEvGgapSHJKfYlmFhgiI/TKenYS
pMWlJMsXW1J19xoR/pyfo1wVwC5VYi+fL9u/GAH4jT5pznbpKqSLBz8wKYbY60c/f0FB8IVMCJiY
epnxP/dbgq6o9BhoJBp213MVIGaUAyNUIXbNchUu8YpFUb15aJXk78z0f4PumHIPYK08riwFYK3K
e/1wqPkvqeF9NGac7gg7dtx4xOF8+NdFHiiMiV9J3neIf6a3RPXpuLvpoqnB3jejUrdazo7wFtmB
la5KIsGIfhfhfbSgqO6wkZn5jBzJiywVl+aGXrLaFxaLMmO4DXSuJypsy4HZP8oTeAqaWdZCKSAx
8xAWZztLE898lLW6WbDeM0GGSJZzCP4hW+IIRceqNC2kJ+JZZ0IG6f7pzgkgC8RtrDOZ7ApQBjIt
sbVGw6sv00Sc9GpwhcXPSyOPkpKPdsjPYGNViNvFRj8UArlzWysYttAhqiN3iXixZnU2ezt+gGov
2P85uCWd62az+6xbuK6b1Km4fkCYQbE0wcc+l4MU5A2zwGWXfydr7lz9avdI7OQzKRy0EYgUaa/K
PsO21abGNIIBQT7Q2YAgsuvEpJb7ZOa0qq4PAPvlcLuxb9kW+afll/pUc9IRpuMBSsWXYC5apPgH
fH/ez7C3q3QqEh2KWJhCZlxppJKy4oMCcLRe0HUzMFEkcxGdlwOtY1dlkUZaDt4CVQextTyr1v4+
7D70wahnNllr/RoeBqOq1OZtU8VUhR2XJEJhQ55rK1aFi7gJjxLtw7ocp7X+lJ7afi90QSIY7sH9
d8IPonUeaWgrTM8K44dAn++4uTxI/H5riM90+HiY1hJBe+5mK0dGzg7QEUzgyfmhZDeZShVXDz2z
K1SHL2OWaU2mABH0VkzJmAi0ibaJrTYRa0hcCYJ7z68R7BDozNIQUkvcF+MTodntP1uhuWAzeyEI
WHq6qSWYNf/dkcZuu29uqaP1OSCFk2kMlFAqhxfgH9vktcurMvbT+33xZan1GSzimt2XRpLKaj7o
fh/7BEYrY0cHEmDDoKZxjT0/Lx3YPXlLoZej2dDEEw6vYv8LP37pER0U2eQPNCePDE+zLwcwbiqU
VZpnkEUi1LjRMGubB0J/HexpMtNH7nQAgUGpsVhNykhFYHBRbLgnW92fpWxqLF/UCGtZIhtvNzp7
v2oqO9/9gRqqCvUSIA1KwpCahYdnIdfLUzltjPQOE1vKhjOuFhjvshhoQTRUVdV7LAdwQKQkMXXh
PN1IUiRXNYjQPLcfdd05htQmqk3+UHtXhJmcjU37hVY0VrgP533CPqaFyLg7OFzsxi5qDCFg4q3Y
oNgzT47v2iRDGPQQWm7VifZC/OMWL6NOmKwtCeizzty07q+k+tTZHIjQTN/WZwO7u3PEztvIY0R9
U7v+M+FmZVQ4+7VQhePR3EUGI1dhX0HEX4dayH9lnaBenBnb1gjONd6GzBJoMCX2rT+YqZyCHMSg
UdZa5P8G7cQypkFB8sim+H88Fv3d9QsgYZRM7nw/JyJlc9UgOEkBuSx8l9S79tRy/Jg1/2gwZi3p
JE/eCPbqcaO3W58UBZeDSJoisVjHdABbcw+O8dtDQS9iu3wZlKQObAgH3owox7rbwdTFyn+WmPKF
QY/BHIvWyGR1FEfJaxOh6sLtxOsaWLVRhEmiPyO2tyGYLnSq4b+qGx6AjLaGkL+LwMGMSaTX3tXI
mhqCx1/DoJDviXhRyrJXJ+80tJoDxcr41J8ouJZ4vj1I9SwzuuPMISwWqs1i7n/gBGpQ1lcjvFL8
i0Po52uhb1Q/DqkcLl5HIrTB2vfg1MsIu4tqKxhDWuur0t4WbagbxCRjvsIN/TvYaNnkC1b0w2WV
/mEAIpF9HZUVN9dinn7fSWIYc46dz5nevQhYR9E/ftzwDqXhYMpDHoCCk3NzEBA7g1C/s++wsQJu
Cs/sMw0Z/NjtUZoU3k6Lj2GSw81wGd093d3K6ozik0/nKipMbyPk2YlZBXcQmgl8jTFI8oF/33Tk
FP5NoYneD8Y0TkVZx8jYoPM79IbYvn4U7NuV3kVbfxT3pVo+c4FSL8RP/8XUl8Jd5RR2G2Cgpwq+
5SDRP+MNs2FapWqpRO/NnPbaOT5aHhi0EbcKwo0Qc6YR2rzdNiL9YkKbQ/9PRiG6/k+PN2fRkZrR
yws5/jL8JEIQNUFIL55ECv6o1jxY6IJYfa8NkWXC2Y33BRA5NZmeGVEAaHGT+L8Z5cTHNyrbn7Vs
E3vLNXUGcGe5dSgvZY3nNzwNY9P4TN0ILOh62U2MK18OdDgkl8hVhesFkl+edwY6BpauG6easbi3
HlltLUmfCCHq2Lvdw01bGco2PFHsp6t3wOAlg202eux5rCrAguwSIdkIQHX7/4dk6OZ0ABkwLCu/
84nAV/AC9lar7xgKfWxsaXX8yoc03Tb4O4ZCf51vL2xC7wTrONCDbMHVkD3Qap5+LwcusYzasnJ3
MSdpk6kpEM3sgWr//rhH3WcAHXxtaZUF4PVyZbpQjl2OXJLIPj8uMxN2GH5lnJCrUArArDZ7VmUC
EbbwCIzJeDKnBXGrIpeGmvhEAxflChI/HddywzS2HjNMqYwzeg2N806R4ZaMMtcdX1SiPVB46ASw
Y8zqjW+7WCdhpvRwLkkC2usOb9fgpb0Kun8w5RifDVxBHuMz6pEdigGDth3U5CCLxme90xK+FXHP
VX9Y/jtMo+WhvA5cHv3FxLaf7ap3Kwb0AbQF24SdfcX76c6TWZq3qV3zXDVJW/O0iF551t7ghcHa
sehLCPIFYkpLq9T0h9mRwoLFLftni2ngJn9B0FXgX8OHvrR3tAiCre3iDIbmxKLZ8JBmKPtJO8hE
8xTaY5QuSHEqqqGs1o/oiviUp9egIPwRjv031UTgr0NuSk06qmq+pCqqzSyNG3RoF9fq1J2/Shy1
ZXDijyTV+kxaGxwLXBoxxjKg1QMfumeDLWGXP71mG8VBtbjYFQUtRJrd786vkc1/8RnetgQh19Qq
hfYntQrCs71WFBmB7s+omD2Zauof+gM1KIvtAjMQ8GsUyt/Xyb5HK5wiN8qAdzGpFnLLgC8mUxTb
3M/StFXECfELMseFBUroraxGNV7RJ0LA4hH2Pv7jGf6nreikw6jqhRswFrrGTQigjx6gakTSKQxe
VIGIQ0bUmKDJ9T7LYLQh481zO3XHVpWfIxZssTOASojGvp5Xb+YPp2Pru3JW72nQ6nMbEjKp4mwi
4TwExg0OcWlk6GJTozfWHEgbf4EDtfw54A35J8FBR/XjSLqYsc+ial95tdfsaiH3NoHut0IGegbx
KGXyNbPpIW32IXBVs2WeyQ3yrfhxk0E/JsWHPsuRSK4YFCXfUgovA75Tnl0Sln+Z0s6pbYf1dK2Q
AneihcgFDXlsS7wRqJgJfxJwsz9Ype/Np0b/bdtDFLDXKr9owbY0e8pEzFYuxAOGomqQUegEupNL
WODMaPVQmvIzFz6e1jrMcSF4mfjBqsUHN3SYNLc0hcZqitY5ku3/bcBaBnfhrQc6aEI7ph6iUMRH
Xbq6IiKNWjRrLU6HWiY2FQ4Hc//j0yegSUZn5h+H/NwP2pMw7U8HJX9cCepiFhj5ZiANuBGCHqK+
z8FXNu6g7i5XbOGJV/oSBaPln/Rkm5gOgUai2pM0OOiQ+cLe/arA7eGYnVjgThE1sBtK+0ltoilM
wlcXrGH5GnaytUO2zCPbIp4iZ9zy9Yi6riMguFiIVTEdGNM7ApDdpSmfZUofMH1JRbXepVKfBIq3
essq8TusIvmbH3zdG4VjzPQse+v3H2Wd2TcNg4t5Oa+TSwUHAcQXlBfOxAqv90gJj07p4Y5XHiYO
5U72uFzZd11uamjfNB8yhRvVKaC70L68Qn5h87Viu6idAvTJAkEZjT4YoXW4MOrsiWeOJftcSmFK
4moAvfRTfkbmpOlRmWDGHJqKz/kQ3bkhfDuTam33CKgfmafd1rjdWa1AOZiCbj3ZEQKBFrtPofgk
KAarY4QENVw02HCpmU+5IYQO1SezFPJsKmQgAw8ug+K74O7yuCXGpB2OU30cSRzuoIjnmEj1Lw4/
8Dy/+PiMZT4XPYK8S9mhRDC037+wxvvuxU3+/rBGRxwAhhvLKZlEDII1B/Bztz8vxC+ZSt+G2FPX
WI3MTikESX7if4tLL+vl+PNrT66iqrpu0LFaHz9/vH2t5h/IG/+5GdmQpyvKrKKYd4+xv/hEE6GG
qu5q0fXi5LAxcpoJ38mUEJxroRimuf8ot0/w4IGPGlgPgjsv69WK9uVWFhoST1+RyXfMKX3hqKoR
CnVM1Yo28P81BRmcHo2gwBRD+xXNxk39JX9dYocneM0TAL5JmwSEgyyEgT+gu3Rv2Q0pDtrckCn8
fdsYCRRXc89i5r6/y70RKayn1wVvpoA6mYdoa3IdDRYuojqzGJnOM7P0sLiGYAoFYlV0T9vBWBaI
PmKslE40ebMcIz84uPJ97XAkb2pZBHdW0rGzwcVyMtz4TGw1oBjzPuMZYt88KBEJUam5sYVhPrwO
3QjxcT65XJHgR1gEeQUC/oaFpUtGfsnhm61kD9/1HIhr7gVlybS+UziFraJBZ2NjLofEHUmkh2O0
Md6DvQPg1SWjOo3ZLiXjgNW08oGynLWnthf2LrVJui0Z0CjZuDbYvYjpzf8n7bSjiaBM8EnaKS6O
6x7qeN2zdMPAmyvoyrWbc5i1lZwwhy4Q0IPd7PpG5SqFfjCs2MV8lCSy1sN27fEwYO/cIDUQKcg3
pVAWRvQ9QLM0mVQkuTzAWK9Jmjq4KfnWG8yOrbO3/ZZtjbzBIYku6dSq/GlhQbmBzpIH48KFF3Dz
F0g4cB04+qeYGxTS7eQtz7I03q1b7VCPYKx3skfFdoOArAxTbEKM6tyJiU+7mffBCwBuwSp0P+77
OatjLEzUiuHOHV/DyWx0hpylPicS935f1ePit384zeawSakh6+N/fBNdy9m41UcNgfFSIreZLhd8
zqpkZGOTFrXpoDG5FWDmP+UsawWbeTrqr8dQcshUC1I6bqJWLnlg5aFWub7ELwkdfpTUTxzYWeYz
7yJ8weCE3LuspvmATjfWxXHpQVa0efmZ5bnVNvq+JLnMY/rbzXlL18jL4yXZ0QJn3sk110MiW0Ir
sq80tcTehXc+5B6/0Rik/61XcryN2+unhdKXMcxAk3XeV7kPZVy43oFl+jcc2S82UWpDJh97LhlU
w5OYPZKUFgniHQ6Eh+nVk2qK61W1s6a6AXic02midp+gQ9ffV2dsbzL0Wfzwz/ykpCkreEqEh8MJ
OvB3/Vm2b7XGTrjsbnCEsoPF0qd+140DX+Zms+jw67+FBFqx6mpuByWbShpL12i7LI1TxFZJKWPP
jkC+tgaZgkYR7pto/QI8sTvh3e3ayUezoEUErHYjP+3lJqhfTCtk8FSz+oEx52Xkex05veYCkzq+
iTmGfmiljGLojKizLVP0Z269TYB04eMw83LLYWn5cuPHXEPvMP3FAtUAnx2W4nCwyNidzScv0CQA
2BFvi/5vzjn4dhM5Fw+BY9syhl1bcw4H6tSvGeri9fzheX8In3FTnXWsjmVDYSxu93y9demT7//W
g3snWzmemrU6jyDKzK1udFip8ACmmNtT70H0z/HH9ygi/wOBkdclbO4aMRPwvpUk179GARUaZl3B
p7OWV3lu3TlyBHCgZm7AQ0+GGxmjYFAMjMJHi/avYz2LBOdgtRkM2g9EebaiPDlss5y4b8N5sMGd
p9/Tu7boz+W/7/W4FNkC7hs/E878ID+FjndHJaI/hOm8tuppAZ3VEBUqwpO11wn/YCx28apWlxuD
7n201o4EacAdXSSkOk+eli+N5i63AO15eh+e2O+AhlXtUfKars5dYYNmIEUaH8uxsjiBXMdX4SpZ
YBxpZMSqwzc7v7AMNYpTWKawP/RQKUllq4+xzS5GiS/JmISkOOvNI/snaO2+b/+tJOnXixhKwR80
HFl+IRtX21zRwmpfwQyS3eJys6jl28Ci0NCqqWSiH9N29/vQ7BECWNNLDXqb7+Aub8T9AGqIDaPR
0K9Mm98r6TVi0MwTm2Ekb8DcobYmDaa6SQt2NpnlFmmkfvDWeLuVx+jfNo7gAriPXnExHGW7GKG4
jC/GBtNk+m8CP7ouUbz64NwxI6YNIZ6UvVRiMZYK41FukDyO8zaIL5guC7mJIP9H2G18bSdjn0CM
iB/+E5pBrJG2Y7PZl/gCX/pY34WDrCmle9N5b/zGQGx6oB6QkJjFKeOlx0owjYmTdk3AJrguiBy6
THuyGohyTfQ9JjcVX+TFbjiGus1vt/TvnR5LTjml0vhqr5yWU33SHE4OJroCpVbwHXU5QX2NphMC
IIXfNX7h/1cyjLjqGkbHdd7WzhGBwE7RZZkls/Sgz9SjQeR44TF7t5EVWOvr5WddaUjt1RUsrdNm
sGde8X52a4NDjv1xaNL1lDzJwUDAIp/v2fsXZJWgsDc/L74GmXDxQ0YHZrjs0Dfh48R+jirpMjlt
tQfk5zoPXIHskJD8xs78+0QHknNcmGyDxp4FCDli7Ak/mqESJmMaJ3u9uwVPvHScAbn8dhVOT8HI
A+KFdq6YAbG/GQfNd3ZxSaggo2UR6w+PVOjR3S0E2dWPIYbOl6VjZFi1YJ7bSjfiE926LAJxiBeO
MyZrI1tgpGueLLOJAaR4aBDI/dEEUrAIalMCihrJ26Snhfv6LjnwLZqut3MFczRUv6UkAQeyebFj
xrFBlbaNsNAsNB4jNdlU76tTTDqFWF97KiLXqIh6tzPhfsefnOfYnSEsbGa9h0BNMRyQDXeuPWw4
60RNJtvQk6+4w6nJX2IDZ1vf9uMGlpvgPNrRxa/fFEg0wFdI4O+giN5Op74M+5RIaJ1d+W/x18HV
RoN1WH5lbS3gFupWV5hxKfWo+cIpJqsZJ5vLlqZLgzZNFLBooV13OOp6VoCZhd13rkpcJ0yezp+Z
zL/Sm5MJeYhnQwO8F4pNm/FrWQAWjbKYqh+1BE3OSimyU+7jUjssDdOps1sFHf6VQ4OqBqrSdmL7
GFNKeGZFMnrLWTG5pp6CEwHhNM82WBbia+CI6qt0vRl3f6wTxJH8e1W4XIUCAc7jRy86fey2vBZJ
2jgh5juHx8PjU4Csej+44IEM+xpK2RGx2L0VoefR+vSLJtGVsgsMqA+yip5Tj+c/sR9HFVdT80qh
NvaY8pQYIUMjhEZ2SY8rm9rb1lazUBf9cu8+bKAX1uswZoeoBO3y2xStjBDF72GOldP+3jhzh84z
DjSom+iKbjimUjG4tpZ1lR8t5P3vla0crLaFxIMVEUW7OGCKQPjT1Icok7HJajtTO0VbyS3+FF2V
TxbLqAmA2lKpv9Vn2Tfhz/SvXphA4gz3cnX0YaxuNodRFkY1nn6mMeSRl9I0+9bsz6QERR1KEgef
w3ztGh/eTsXkufehaRRtnbHRQDCdgUiLZAT8BbkuYzBjenn9nlI1Yfyu+TNBf7P+GtTvhye3Vr6Q
OlKyA1iRb+X1amiywmmfh0RNTik6vVJr4IpB+XdpyOg+YuX+JoOt5bPz+iYgaAy8vaijz6E0S+n8
Gjm/CPAugLuwl7BEbqqmydDF4owXvfQO0ibSUHPWpLgv6yCRVK3mqMvJO+wJ4ykyjIU3+xFg2PKb
6Gy8WjAWGMoLLfbU+m3EhQ7GOp56P5nHjebjup7JpOX+UiPULyie9gOHvXmZak6NOavFFQZCw3ZP
lAlufddtyfSBi74+Z3z28qFLuqSKaqbNtxn/VNh/IrbI1mp6VO/61qXmgBJizXTse4Xl0+JD/LMC
qcddRJCnn+NFmtxWOTyNzHowACSiZM2UNyKVRwRAf8VHQL0cJPK9LkJhtdk5pg3YvTFBnG28GDui
IuTumaNfgx/Qcq0ZWNCV5hHJnI/HDqINxSDzbh3Xv9ZOk5sGrvmHB++5yferz4yC204uQnpyuXbq
I+BuEgkDamu5yQ5znCwUV1pznmFt4cNRJS+MD0GURvxbBInTWZkbej9J7q/cOCzoHf7rm+pUgjYZ
mc57GDUod8kSjbTKpoCbJrbPlyo+a93Rg53vWULWZcXlFtCkXAmMlSrMLUOMXsJ/ySziRo2ArZlx
pPzPUNQZsHi35HlyPXXDnGGSWDaIjcqvT9s5qamkES3b1aImCcsQWsDph5f5GtTGnbQ4OUEc6Z77
5lXmdYnU85esojz/PCB2X/GHUGt5dbyd++JMWvyvkkyDLpQsIq4KFCGPlT6WafnB32aVbPJ6Qe1r
r1p33agTwq09a4SvKLKdt0G3KCoNgdPZgr5HhApeC3NzAIlE+EKPAvA5+zsJ/j/ZTfPZKde6wsN8
Kjq8RhK+O9ibq60wWKoQ11SLDplzyKIrKdI0kI/RHP7NC7WaR3Q8ynCJnhfsj27z7DPoq7Yr+Mhi
ZEM/7mmDIzR8JEl+1OzIvatruOdoi1AZTktelRzBKU836vyOfgQpAv4X7NF8k6W6up3Bmw0CwhR0
nT+T8IC/KxFRIW+EGU+G/auPFRjEM/T26ztKTHqD/fO5FBS/dLnHjC/WWX0UbJ/sn4koTb7rsJlC
J3ThPThOGJvTfi1NXYkMES8iFybijkWApgawL47YxBIUXXUyBD4nPZSCvGvpCFN/vPbDhOICa0ml
r0RmuE2jhOe6y0ULbsjLxH7a5t3lYUAll3c2bnReDDfXNbHZJFfoLQJEf94uWkPSsvO98D8TFsYh
B6ZrWaPIc0Ikz7bA/xYSZbaqBoYi84v5liMTs63uzXEzwrSBEyDo9UhiT+4FH9mRFKvu2enLNMU2
UsfXD8w6WlHuKBWf0Msxoi16SFBXRP9NH2GOBvJPgADCzZQVc7TK8iRK5SZVoOvdTDcf/FP5nQd3
dLz+JuU7ErPeRw5G4hDWyjY46ReIRmTrVXXCHtSltj9mtiBCKQqwebDpdcm8WkoKLUHvuss2W1wa
0pXLmEOz8o+ZSHluJADqIXVFkKdaKtp/ZgOlDlXRi5kLEp1pXpWa0n83BVO3Rt2JWATa438GmHWE
AVzlPnbkFgE01AMI0uZ7E/17QRKVFhMhgOq0jmTGGsD2kKwpfLstZJg/gcXr9X54g8fGUauSx+LV
1TiWo/d7anhKlrb1Syq757E3JdpvBvPVODxpa6C1M0zeR4L35DzqwHgYxIUHw43kLw/jpykGwuiw
H/7dYuQbk0sfo0daNAcrcp076PsQxsj0Ow7tPGqn3XfQ1bMGshvepktSJixynEcb5Aqnvs3s3zfT
VI+weahKTjMYMmFb3Z6KEwLifby0/pCNFni3gs3NyZZK8KENhHMowx0+XcK5TlEmJhjXKg5HcpK/
1k6AQuobVWmJvZLtip5+A2TVZTvtzxz7dMSbk8QaxlfgXmKCDDz8In7tYh4Xra49kl9wGM38ufiO
hesH2fA/fnryoaQEnZUqtl5a2cIwlEBoCRDU9TrKQ4s1Aiv02V2vZz7LTr8B3QAt7kifFqG0q06e
e9UjXLmRBDqNEmfMCdLjATcj1lebtDdKBtyhVaVNJ+g6Rmky596fkYtMPOc294ncfRlhAtuCLf57
Xf+DC7Nr1bXi2Nl4fEi5hsvkDlNOFzpPEuOU8nzXfYXxHjcg6CHGc0IJcOdSAReUxIS4jlmW3GJc
QmQxwwN1cpt9+zsNgiuts8eTVWpdZ9y7OGWWs7eM40iqikNFaHtc6Ceimh4NbSMcIp9r2slW2oJ4
na2GaZKWi/NOFJsz9PLOXmzP/HGlgt1rHmxu5/d42hB+u7HXCDpyE7sc3bHsQ/2jtqDFBRNsdH95
XHovONvuxd69+y41KeasKF3unB6umSGv2tp8JDtqr3KS905vEsq4aQmhwK/9SQJav/6PVUlKrt+f
b+cSSUcLImFYEaqVL+fLsQc+IQee77inuIyvYhRl5/OGn8dFgEbAe8zIUAYgVbQnfGs4Bq0dWrpC
nzFHz19mOmuAHjnGawxcLt/Z0YlcVYnjBZZD2yESleXlCoL3KDd9hhsN22ejUxu+2Xt+TrkgM/HT
b03/BePOXZ1PVNXn6B1xEsO8QkWjSArzXH4vYO+1fLdhXRRfXRnTaML8i38j8qEbZMXDHM7fqYRY
BNI6biucSHa7J/m5zB6LDF5gxNshkCWXXwov5HCNY7HwZ9vMlh3Dm5vA9bii8aCnxOHWZ/zdykiX
0C6SpSoaRlsQOhdeYkYSMND6wOGXOpNceJC6EzLtN/Rx2M6NW8h4tnS0HYW2k4798wsxDArhqSUd
AMaFVmMBjlpbBmegyk55kSu/bEu+2uqaOMGvEuv4Pbx7vj6MmBghW7ATf9jkkUxg1o5pr+b2Qm1J
Ip8ZWbE/JrUnbwRKyyns5MS+fub3ZBTZoIkKlNgfYGkK+TDwBRihhCXj9K4/VF685rzva/3orC+E
pIq/QxEmeKuR227Tsw+SQrniKlvNQzNexNsdx+S0JgVQTXv5WDpgoJp9l7BBhuQavscNo1km/t1H
LA3ZWG6bNSJMGu31BrOAccpYyjMLYkG4k7YJO2GJzxdvCLbQxZVb7/+iVAcZp9WerBO/Nt12t7l4
KdtSNkDMnpB1AaMw+N44wvk44qVrE3VbJZ/b3LmgjSQUVlREfBNJ3p30KVybE3KSvSJgLyi3aeGf
+KZ8qHbrQUzrYf6to7cTLrMMiwFe9zNNfOeAO0pRmysXZRh8PmyO08WrB2PGO8aWEPd1O6Xj+Sgc
d/m8kvlwdVPRyNYTn4iNOFvUyYMGtUDfK0BNvJQUr7EpaV5sBNDPjyGiyc5LZZmDLagbO2twG5Re
KwOW3I214t6p2Mvv4Gc0raKbZuDEXqL5ekxx44caGuI2NS61Gn/Dt+IQ8ytfx6w/uwhTkxJkp7IY
+jhLTNyLKhIWmk3w1GQgO+VANAKjNFb3RKEMt3iAgrotF05tEjyISF/JqShrtVlJGynLnaKOcYYz
Jxq85T1so3Q05Ct9LdLnejiyuTazvsWw0ZfTIwsNgpPk96H8GmbYc/oQf3OOOOB3Chin1k1qLha+
c5T+IXU+ny5YHorw6eGJtBkLfRScsTueONvld7F+fwEUjH5xromxXvY2Mrhm+asQZX/f7YV6Hvrl
lMEgqXGqmJaesjQ7r9B4BdjltkO5j5Qi2tRDqgNGmT2W9BNDAoQoQM51nqZJBkCNUSZ8goLrfyAc
ctNOJR72s4FVa7zO1LdSYFyn0WyCCHs1xJR+w0XN0hkiJJJoU/uEA3uhd7KZSgiHZx0h7QE9ZQeR
dpMxyZ6B+0e3B0vtxBmXAgFygIPN5zat8JA8OwR5t8XYON0LEccj2WgcTA631zOJI7ERd+8XRMhG
cYgeR4X+/wpRaF0nilvv0iadf7FxDAUjHGrOFJYUhhtaHQoHqDcZDu4gaNMos6adubUk0H/tHjOF
AJ9Xr6J0AmYC65O2ul/caujGsOB5Qs6tJ+OvUYG0dCGh90kkMG6Sw0czGngHxq7KZtHVhoW6IXBq
UqIDeCdRcix5/C1WDfvRtQKr+wwOWmF8/rwdA4GqNuE5bWbMtMweyRF0bOVbXD1d9rDrE1VopyB9
s+SEMc44y7sO/0JJ2jz2e336xQw0TD+PGni5LFyvGNzkNrcrHqMGv5L7+gRZ0EfMkVcgM2plBZpH
wtEsEkFVIkduwXfR9X7b/RAFUawm5b/bnIPxGGeP1XV29HlA/CwIYD/PwfTU/HxAh2in8CrqGtZG
EVclyzQFQ1J+pTWBWQgOuFUMSLVolTU+MNtrLseu5gYRtRVLx2Gz5qTv6qkjZjcLAilQFbxFsC+V
LLZ/DarogXZ4H8fDYcTlo3s38UNXtTJe9gBNrMqh1m+4yWgxL1+Lf4un/GEwf0YUlLGrAx4nGlAo
8kXKEyf5ZCbojAp09/8pB+fAcXmlGBrp6LXmAg6wGWtRYWSaPzypOAYWY3Wq894f3f7hbRDusGNl
VXzSWoiCx8pb2LJkFimFmmneuaDU9JB9FgWyzc+Ha3nO8E06BUtFHLLKZbs/0idmmCyl+9LDiThK
rm/95D7SctdWIuY23WCXuOk9menPeZNLmes+0vH38iyVuggIeFWQnnejI3kh4ZLm7e4NVHHMjxXA
DddC7beGLq+3U8QhngwbUYiu02NJYC7VmVUV5+2sHdcCaC0M6JCOAQdLTujevs0MQv2Ro51ppJy7
iUKN3uxl/Sd8k6nvKjvwsktSqGZO6AJjD1MwADKL8gvd4Kt/a+jlxncbSupRLnP63nz9rOHCspn3
doNm9Ka1rXg+0rzBaGs9iqFNIVAxPguWfpY99uhgvNo8uhuIZgGonVYg4+EldUFnXOsBvFC/BvB7
g/ZuWkHuq8StOMMkSBwdU5hIMTrATK/dp0lBgWH8T9TNkFJJ86U7mVIKFU1TLLkVu5GXBy0K3JOJ
/ecgSvi81BjotMPBiR2/KQ+aSagXZZV0ZKxzUctXCWydKg1B2bX5D/0+YiwV50NNMm7JjQ5OoDt+
on846rO0l8PfeauAn19fK0NkF5oOKFBsfQYOQpwWAzexuBFnnS6wS7QVQ1moHMSUuhxo7m0x2v+h
J7lV206F24y9nzaFAhnSbVD+XxRepdc5LKtstZrBFfOU17pcKeAw4pecVMKP1d3O5AKgj0BEMNJI
f9dKjo+g7HKDK04P+u48zhYQvasVBa9mDXWgCj6ok33LWyi4KcPDZx5OdZYXX/oRnXnPIyGFN8bc
ydpCHMIo457ikPcH4JTTT2bHo6Y2iCysAKNFEbYo6dHLilyYXTxr6Z+orF8keDLYWQGnqElVAuRo
E2/ftqLeDj6H5tYCSor2UtpAzfP6XdIe5l1KsuTvB7j6ULsEwsiZrU/97iBar5Dt9p+aeUvUgNr3
xPiGNNG5kJWCUBaBf5p9gaylbNeRzX9fFfT5g/OG2/RPgzOKs78Sik7G9jOMBReY6k/+B7JxHMlU
+pq5mdQXZvMz1fDGqL6hWzsPxHkUh7oE23Y/IE/VZ29clvdSRDhrSS84ehNCLadmSrdJvBpbOMtx
se2gr4yH8HyTLGTDFiuf6MvdBaqtXG4H5QDP1fkznG0C01gLF0eOJnV1Bcyje3ru8d9dLI/KjD5V
C8j8vF5eAsOCWBd3c3cALn1QiMT+dWk6mMgKBuR2shq+IuNjCfH6u8LcMyQ0s7bNYL3vw8h9szTk
EUAtFyYyIEo6a/eWeEVVy3N/IMvw90ejwk3Lq8V31MH/TPMEi/zSM32fPKMfTNntPkXISB/W7rmS
boudQN6ydNWp22DpmbWx3EO1Wh2rq2D4vVscFDmse6t3AKi9lTA+Eb547htK7ZCoc+0mYVYURv+p
S3zMdwq1EjIm4FFHo4kN/tDbQqXNvpRNY2/7sfr64sZ7KWc7x4ckjgwusBOaX7iiqUmXID+8pRQl
RFCJkmNjo0bhxhruQMXSnEg4piihSYnpY4kG1NLdTh80YdbAsq5y9J9yefg/tfpslJiQHWMb0qgX
22DgRkfz5N/hpllFGPEOZoeW79itCc5lWQbcE55tKO2wOSQFnThEJ+a0ItMCfHpf3eNBeiUisZG6
gvlhay21UJS6xli5o6HGBWfS1DW7gt1W0wLYj0PNVtFJC7T5CzaKXY/q9onC/dUKO2Wejl52jjPf
9hB73lBFyLqwAYEJJr48KlMKPg+bZzyf6xVRYW/QgGTxXwsvjXJMUvwd8M2wSWakME26rYfhYeIA
hHFfWD2yAhbucPtpWs3YMiARay5LLmLYuN9JVl+JdhQWhyh3UZWuc4INyQST48PJUjW0+sg8s8ja
ZadRD7MA/U30tfnA7AqGZqf/QjFRZrQTnwtaxVNi0eY/mmdc2lkJcUpr0cO1NSqtyg7MRBjZjv9k
buHDUF2ux5Ywd/8uDHQbSzrdpO9Qhte2UIW2t2xgrmwinbW0HgNTehia3breFBvojpUyQHKeaHA8
bAEnKetOwgKC5tsvHrmXl8GuvZGMaSP0jDD29WebU1KkMsiek76rz9q37nbJf11wj4IwJKxloL4B
ehSAo8yT8V43dJFH4xVcB9s2CoEUFVgtnR2+q58/SvelvCeUa+WQn3V/4WopLZMDN2J2OadROk+g
3nfKRHmGy5VfPYeSK9ZNmHPdykB/wFYNBuKSX2nIkwtHM821GYjIvgfHUXhmkTwy4iUykPxVQtXO
Zq+FASs5f1ekZvDffQJWfkVK+ReGQOgACi0P2oBl2OREq2dHWcbx5UFl2A9wT9eo208/qAeP3NO9
0I97f2gFV54FND9RCTCgDoRcKjxhDAwSAyT56F+M8uFbyZed9InkdqwwLrlVhFDrEXU4momt/GIG
K2ot7dwzcwxOdmEP+5jyTd5acWNG7rkShlgGRxhtHDc9gGocwoGe6lj6cvoNIsSsO5sbK+s9YN5H
Z7Z8jy3+ivwzyZVJHThqwnBdmw3ffWX9F+CFNaf9UDJHURcOeXpLn4GhYppFNebWoQhjKVfA9keW
ExnN3/WWWzOk3oRdtdORXIkmrr/p6eifSF5vTtbW4krxMfw5Gih93qOiDk27K1GZRBQ7JfAqzoFm
5DKJGH3EZkaT3aMOA35aEvi2ZeHtKhwea4jnkcJ/awRf/zwprRIj27HEL5kVnNIQq8FbhtjYShDp
r3A3FW9pTTYNuZOaVYnL0j0z/9aGyHSP8B3bnQs3IjPNyukI8AyQ72uWx9Z0W6UZZSXGH3BWgtzC
zcp/EudArInOPaXbFlyj3RHDV/688j4q11QU9DfV50a/FvbxLA02l3B8G6oyTlSZ8v5C7StbI8Ls
ZqpCCI0VBGhD9M5ZnBQWavxK4XExayKQvjPZcqVsLpYf4R2nzeW+Sy7V8SpLzHeL/BhHedxFePuY
1rvZYt/wi5n3mzHXWxGs26K65Gjo32esqAV2cl70oTBVZVTpvtjvBcuXyD8GuQpD4s8nNBh4ywA+
KS9+lQ3IVqm8gxLWG7jZiYQlNYv9n0L9YgDxQrNtZf3VbrrogbYKEQeGmy7pF6xrBAWpG+2EURzl
JYxEPwwareulYQIa7cnXLdU9PP40/AeqOX0s81GeHAmiDGkmR7fkG6erBZcfgy09zzkSvHyTUgsA
tqEaQgB6GQARTB+P3ol1Jc+sAWmkyeprq5/gT4XGZi9uaKDy59RQJnEXhE/G3MNcpCINBv18SdPO
WXWGfAdTHBifEDOVmYoAvJLqrylMsBQH9MQVAhcR7K0oBHCZ4DJh9MAGBAxKH2sR3NXAGGDlYBcD
prwzbTTm8MIunxWUZjwhPNdcUEepm++7CMeZ+CJjEkcj+f550w4RysUhOeCRoPYQbzFlj74+seAP
lhVl8O7S2wwwoOSYUkCAfEb5yZuMkhRO+QGfvb9vCsQUnpVCHkFsQG5K+6egejZlywkNhBZKBz5M
YtnBqIKcmnCpXe+fDNPaD3u8ApecKjtp1/uEk80R8Ttf2MfvqmGPfXjIoII5kKXZFiwmgEGOa16v
gcgItKOtYEDSU5qjIzj47tjcau3a/Hy/4QnJ6coyhIO5GL8WMyJ1PQC6dj26VfLbZgCIfJZspmgE
DBUeORPAiWE+qJkLJ2QLLJ6csXdHzvVconjoIN6tsLID1ZVX88mWz0DOjcBWxcELa9t3w73EMT2R
sCI84cJPF/bHkBrtQiCUkf/1TNb+yDKNBAzcUsMm+5wKNyRaMGpIDR0Bqcv6Jv7aysWDYmpCWfwe
+WR6nEpm0XykFir94NBYAPNmQQW6JaX8EmmVglgWXsxTOi7tG+KTIXY7JmZsquawJB0jMrjFUz0d
EkpZoz8D1BrJiy76F4MJDxpdCvgpDjVKVQKyYeEBdDgZqYL8PMSCfaRUhHLKfbeh8M2HKKawzzPc
93sSocrD9m+W5B4CaFYh1FPTIT+2KMdJgJ2r7pgcP1/WsLqYf7/QZb1xoSUxHGhcCMBPO2csHOSV
MWYEA72P2/NLGG+NYqcpFIC23VLXWKAzilBSefibza52oz07amnHRMlK/Ac55qOHPbEJo614IPEv
n3SYKj80gxpZdngABhyKmt3yCYrclgXdRfWh4sGqeCs/O4IEeFSmCsdt9Ijfw3Mq7QyNO7AIVs/s
L4F8NCEBSUT8yA7pCsjOPoTzY0/broMag8rue16f5e20eU1JCyf0uSnxJHSYD7QMVcPazcIBNFgj
fUAPGQn9u0rU6xOBn/Qml/CO+gsZUNgIq5y51hHrGoaxCXJDG2/f5kWMx188TkQuaqRxCMfHTR71
OQlVsKyfirxuqy7NBLFUagHq+eAJl0rvKOjq5P+NxKFxi88jFKw8kZgTKkZJp+wOujfrPIP0go3Y
all/G/sFr5Lq1iizorWXLiw40su1U5XTKnsAF5euGUUll4TSB+3oe/YiWyZEUyYkTPjNiwQFcDaS
OQJqTKzsl3gHT4v5vFm2cCLaCVeTJGFrB6gITgQHy8m/u3FWhn0YlN1+Hj1vUoJE2gM4S6IoIroi
Ee/xWAtyos+IdY7LsThml/fZO9tV9xTHYFZ86GXPfoI9onc4yGLsEQSNjg7KFZe+QvBlrYe/RBWv
29D3Tjxagz81ko2UoJmjtfx78Wit6dn+sbz7dS/p5Y7WcF0Teu/FVkqzTNTmUj1TEHGzLyQYccw5
HyvEuGkWfJzUKdVDGsgi07jHiVVqduyx1qYD9ifQW6mr2wxMeh6yu9FNPxO+u0EbGECZV4m9D1AQ
VqWS/cHd9kasOl9/mB+ojAeJhJ3O9E1GLJirjUNRYuUIEHG/KvBhvtN/mVPwdWt8drXHDAuXa4Ky
TSt+1hsjbS2U3Cf98qhPBxNXfbZBffoffIJhe6OGhGYHQ1KPAsxI0ccukOseWbW4cbrAqgAJ1q6Y
sQc6Zqh/+0qO4cOca9m0UPy+r8G0Sz/Ux4NyUFoxxo+shbge3la1txbon9fx9zJErsu4f5M5eJ71
qi1vCEsTb70ves5ODn5u9CQ7TrAhWQ4dm17RePLyhU0yXNXgxp5HPxOsx024CyHn5JWmnEKttnAQ
ijfykhxd8bQxMTmr5mfw8hl47Jc2BbTQf3nNw5AkDSyrdvMwXn9mXv97GEgrnq990/Ju/lLjBfOE
t4nGXGr35Ox16kH5KN3C6G1PzueqyLhumiIuwzCAG6WxErQOyVAPvivkC8jDWFBiLYrRlGgUanS9
MBkhYIhNJpoBIX4WyBHsz5VZ5HMF2j0+zWicAqA7yeJ46vxqyoeMZ/QnkMrIWm5SNgOAVAIs0lYy
t6W5mLy3Kcp5REcxczSktYT9RLUyA+tdn0mobhc6hjnq++2kRvNLn2G+C++UY6bamut/Dim59NbL
ViAdBdy5VAo+Zf4qB3GoWhp4BKIVugwRM+NmnRmgEt1xQdrOC2OHgtQfLNA3VqQqCXGcdMeQvIm6
ZzVt328x6Fz/j7vd5hxZjyB++eBfNQ4Zk1QISGUxKsiZBrvmXyUhu5rYf1ESrnpcP8H7pWoDQqPb
NpB+q8SaU0OXkQSHvL/Hp812KGekcxSsKAk49hkrlNsdnd/qIB0vS6CpxawtrPbCiKdgELfKTJkq
IQ8qxi23Bhj1stew+fbFq6jRotuxr81dZwQjLMh6PThr7CXsgMgzoVjoHAvGN6M3ioZ1/WNNC6Vy
jlrtec0W2GZ6aNjeMPUrFgipLQvt99Oo6377sIBdDJGX7RkUtkhlPyrd61D9ZTXzhKXoEmlVOBfu
DF6YYtef80KFEKodcOAWvx0rzn9Em6KYC1Ley4CeEhf8y9WOjmI7MYQV48vw+FIlYAB62eYt1iDx
bbMg5VeEmHbbAILbIjxGnH/rr7ZA5KKedr+y1Hzykp6gAhtJbSn0WC6sjK2jJGxceBbKJgeDmtiH
Tzzt5wP+2Kc2wWoarnD9QK4oTZrWmUA6prWjN81efXkTKs4MKCqTQwQONHj/msSeOXfYvYRYStm/
yZkkp4/UaLDYbmS3d8Tat8gDxhxsbKoHHloRm5A9z4ncSFwwMaexQ+7JAsdT8bptMhSQJjsAkVp1
QnQ/e4s8jcOg8Fa80MT0udHFxKuv9OjVwL30MSMsY5Tia0dSOC2ZytKdgGoKLr5kyb/xFx5noTms
paH4ClKC0S22jEsDLeqaGS7j4eWC037jenGEuDXvXV+a8ut2ZIaq/Y9EXzsN/b6RTmdnWbs34s3D
kB3si24uhPQvGUI1hakCz4e159ktiHwREnJbDpqecqZMGrrtBO1stOymNt8ssab8Yi61Hgin9GDB
g8Rlw6V8ElOdqzkl+hKXge2AxppzFLhfV1WuvYWidi9uKdeCb7+2f+sqQarK9H2Dwz5ikCSsH5LR
JQ3AkXbCZydRC5CEwNh7r7fIPn+5Q04dzU4EOKfFkTe2cblM/UPWSCfDTP8wXbCUgdSuPFHj8oAX
cr6r6/XAYtwP08UCwNOjJmZQDpoqCMlWvUNPldIsm5SlKSYzO0AdqRrD3XQ+6djSlJlVD+xuiLHn
Y+s/vHoD+YfQ6PlaQ1uZwLbKy8yLcGiCh5rL8ptdFcrvEFjhKfowHl2sR2XzaRlFPV6S9C7Ft2Sk
YTdDMF48rv6qS0y/hwuWlY/cMu5OmkWN4yfJrfjprg4Cja6vOEkaWpoykRp2Mc16g9X6S633peiI
tsTB3B8lehSXiEP+tMXWLSimjuwVyjyD5XFVYVNhJuuzNNemwd9GS4Qt558B9quvCL/EpxQ5ttbL
gaAcEx4ZW4GgkFVG5VE/D43qhi6adKJ5M5WLh5NmxJfgGhSWQ6MY1IWJ3CSTxenS3nqQR5Z2tGmK
06mX9nvT9JwnLcbqr9IxFlh03gwYRfQHTJoyf00KiCTp2aZGlKMTx7AJdAuMz/Y36aUfHFpEP7kn
dApHG0ex7QbF6ixvvQ08BM5dn8lIfE7lHkhTEhValwrRNslFekg90tjfZrNmdlH0sNwHRESmTNZi
zaWu19JawHawkGfo4vUMO9AGf/qNEgsv/kkwEBa5puJa0sCLaKPZaSMJDZjPlHwaEAaY8zU8/5ow
n/T5uMEl++afyosnZhVMLzrFgAXPUfsiekw4fvz5Wfnc9OtV8iQdetNhmaBMHhZnhNzyVjq0Ttzo
zn7p7xmh1hu/c+wWmhgweNiJcvOJfUnISbCQZS4/n7wDpCRWW3szLRl4TI/wJ1UiO5PtyEZafIrz
OOdCEjBlarWIQhDZEIRxtlCmXwT7a6PO8aqskfDdb1BD2UBRiKPfaSO36vUxVqK3MGUm8h/g/SbQ
vyAKbn980KAf4FF5LOjcyoR4TLKYjqNkxFqimeVmbptl5QjX2pJgH+oLSVBN+q79LymQz3J7c7b7
TtgabmKLwv7/YP0Yjvpt+RlsQVpRsKL2haF8TBzFlBVZLk17+tOhi9xX//MjPtjbr6WAGMjztcWw
t41RjMkP3ZHHS8o7OaHjc4HxMwSAQpGHu25EqV908sg+DzAste6xQEA6sM1bzuD/V5g/GGCyS7+2
wdgKT3cx+/VLwYSFaURw7mt/d5i8Alsgunadyx8NxyUdVA02nma/ksxccbhzI/cAi+h8EYaCGUxC
5zh2TmHPgLYetSRH6aGZN5CEGIlugFdQS3lDqZQxZQusclFtb1EZtsC2bw+h31gCuR8pAnCxfMtd
qk/nQOzdyIeCEPxmcNyx4SoGqdofgYf1VY1mpKAbDnw3LUntTWw4VvqMekp6smI9R00MAfT/xA+u
cp7EsSkszYmi/6Nq/2HeCVJ87i99L66D46LGDNB+TvSRms2e1E5VxLAxAgINDWsH7FTAfwLuhy+I
LpT80mGeqdeY0ORtq5S8xOXeYCIlOPiPgchgTTAzcMyXG0C2/yRguNqauI6qKqeJW8qhCB4WFh0+
LzWgcAn627eK2QTTqk27e07Uxb5MaFoQVPKihEd/QcfzHwRQBC0FpInjWh935XSGrj40fCR/Q3Cs
lOOy2fGn9Qh2VGYfLfX9LMoDizTBP7Y523iV7EyD53QM92L5imLI/nIqoIw0mH2Kn3SToSCsGXe8
Yi8hC9GNbx2PN9tJPukCI2l4YDFLmlqZQChSulyqAuUbCzNe982rJveX+SzMOlpq0Pyy8V4pjgoz
dzYtpsGiVHMX5l3NJ816zM5wg4Cgbl/xmWZqK7uvwMaoBi0wxGKg6NrDxjmX45WHq61+nM17rtKL
gW6UD+9vsOT1Mh1490NsObHHQbI7JoxfOStLhbZ7bW9Z/Om6HlGeqn/EbSoD8AAXEQWQSWOZ7EKo
SkWuWHGoddw1NS691URmw2JwllUcTxZ+1vm6pQxoqffrcuv36aZ4KurCdvz8C4EKEvIEEhgfTTCi
dg9CGBNBRp2WmA1V43nWSKcpWqLbaKtpZqs4bucSWU0//sNgDVshouBksqy/EyKZZhSRXbbBDieg
LxyyIurYxRry5rd5ecHH92OLhMrW/Z0KwffsUojD3lEDjFfW/Ddb61VhfKPy8FL23BKu1C0yre+l
vrn0hL4b1JUcX9DHESeS21kcxrZuzH2cDmxdT6lTazLu7bratea2pxZLOI0hSPw8rd9A26A473xZ
lX0XS5zPilAv6j3fUcZF2Hr/UnHiu4dDvP+Xfb3yzxiVxlETUXrYPzk64X5ws9GhRzXZqaqG5vdo
LA4PLQptRWd/HvzKAietobkcPZsskOJFZNg40CeAnzfHhFwxKk+iZYZH8B0uyPMSxzV56+JMGalG
TfBthe0OAR4/uhLYsZ9dGfLfIuex4cqy5JEd6LtbULiuXvdl2C/MmD3FC6b92yMBJpBMlcm7r2uH
dtfbYZ1aIZTyuAQeKHtSsydsotYA/+HDcZirWs8veBI9fZVpfLJZZUOp6+nU7Ui4tzZ/bkF1SdV+
3pjeRJ7xsFjWCn4956vihAbeYGKmwX1DKyhq9BFRGif5NZB/1g7slO5Cz24/RYznJnD8Nr6VMnwA
0RIBilqkPb7sHBFuWeEXs57jnRX0fJPEWe9E26+kUYGI6gb4ie8QfV2W2/BAxRbUnYxu0rzUzzVF
LOX5cbTMluNzAeh4FDgrwyoQVcCh6Cu1jjzlJL66Zp0k9Hgcr5VoBx8C7v0zDemCCWTMNe3eJExz
ZKqMtCDxY1EoIHUQWs0hIHDdOrda5BVQAMQYWMmR8cprpl6WW6/svyRiycXrmiK4cd32TeZM/mcM
IcTaKbWeVw0pYwRTwgZ0baCdpCuMl7Ityi2IlJf0Bv5ejZzt0+z//eBNaLpvt9gRRwTOagkImv+5
y/Ncb1Y9/9YBQpxVl/HMrGyHH2U1DbpSdZgO3zEOLsYqOnrWxSJe24nOUr6R47J22py8c2whleTf
5FqCtoy1IUHACoSGzR4/pPaxEJ2L1E+HxMtix22tYLosBHpIu/JqTN83vFggWC19l1BwbXF/Y5qt
y73NXJfstnzoXlG0ApiAzu4/X7w73cPUp/D+SQwMIgtuHbLIl7G7i3QUOoUHdysg0162mH/nYa1M
roxxtUFpolAotTHVFbWzFhzbXTlLGRXELiwcTEbYN8i3cgkWQYsgaDpr5rGh+pNhoWJzfTZ7LnWy
a8zJKarm5ZFpkqf40flwsSjyy/qhz3NT5l2Xem5b6YyxxTYGXJY4uwUFYu6qAE2OrggpkzRm2YHv
z1mOyw6iubbOJJuScYRHk1vargg1nfNS3EijqicyRMZ5Zfyz4K+KiJ5A4cQC+WUL7KeA1BVf2hH8
wV74bWxNt76R2D7yocJiutJD6KAEqIyNR86zFbAjdKDpY59kV3kubHI2LKxyPIOPzXwz1biq3m4d
sSbt1KCL5i86qAVuIqV1cT0jiJ7onwj93nSVVoGIeGQ3jqg0QGlkb7haIw80SujX0U+iolV0m5gK
BbKAbWQT65ZBFlfYH4aHAm80E+yvDhJMx4PiMVyqmTUqUPD+KOT8P/HjtP7OEVu+7WbEK1X2q9/g
vFlvgw/rkSkEVrvtErXs1QgYo1v5UNjszk9EyiUT/qVHBLkNkXbUJJr/4ULSDGPXxYk+1XZZOvHf
Qbbne1P5AVyprtUyX/pruA/Hzv3VePyeAKtZNFlv8vjQojXIlt8nJDKBv4xciPVl04af/6qQ8gs7
9sVoaKpvWIaVoNoBPheM8rQfWHFrrhMqfIq2P85Va775m49ZJi/AQyA5Xk9YRl61WOig7Wvgr9bL
cjZ8RrtlCHqmgHnvAo0oTe+29lFlp+MBGwohI80sFNpK63tXqHsW3W2itcPoIs1PZZXU3/5tSSIj
Xh7JdzkvD4QqBaDnr51oOWrmj5SkEVoSyTIgbnCq9MFGCX/2h5CBJP/JTFIwi3UG1EO6lWn+jcx9
pQik4gFkZS5cN11zyir9FSOwVkbhfljjNRG8GINJJLoPhX7YdYPgRV3wuR6lV5KcBDc+zsZdYEJe
vJqACzc4b67cbA13G6WX2U4nocWx6deWGnA8VmyBdqwmJc0la4Vz4UmocHCAZQXBCg2TStFvv4Hk
K5K+f/UxnN4GfzI2R9pU4zFKqzeGAZb7CUDF8UCv9MJ6OFDiLlYY5FpkOfIlqRAhbL0nhrHIAzBI
PYyAa2kk4H7rwnkquGey/0do2hyS8L/bKArhPbAB+eL8HzMJWJzP7OWrUJ2Ht443O/ZnGN56Pdxs
cQbVIAQKmV6usU6NS0OCGFrZDX5CFuwDtFwJzRDpVmdAAxkABUf2gH+TbBt14aXHvt1Xr6VBw/PF
lm+cIIYdjOH4ZL/ftsfyBIbuqwzt/wPIMmWXkl7pSN/a7AvAxkX2N3HA3sm/Ldyo6w07MDrzh9KZ
EYE0AsSUkB288r8YR8Zsrr1AsXDbs0mKIqgPbw67b8+ZI2OHVijaZR1z41GFqT2iBNkJ3IWMIbI3
TaFMBdOxkFyYqImstTU/yriwI9cHDP8+fnEhUuVQLztpkIoSSsntsba9mc53kt9V65MZGLgdeI6b
EmrojIseK8YI3i1PHBXf0JoCRRk+bTz2YVTwly2Qp5NyoY7hAEdIH7iQk4PX9k/C3A+YFY7Mv2sG
ElSWEzQRB5YuAROBzrouzehutt+Dvu7ugayQoRnw6ffO534DdG+CsrhOD8NKuwWcPPrmequiXyoE
doZcafOOCweWMfuQAJnpEyP15Xx7/VuAjAPHZ6OxmAMhWMEiAH3UsSxUtUXMEm7DohPs6F84MYgL
BbwmkQRcnGQAKC9cMZdq1OhZFHRrWDgfASxfjRPUAzPNX9jZDDBm6zQHKP82/WP3Z6kZOG7cjyA7
KYurV1BrXaqlCbsee50ljNZQ/iN3+8sRvkvffY98USymUFw0PNsYhYv0fhQI3TXBeCmlqYqxrxyz
tq+aInUYwHZs4chHu4AvpqBMUtJcB/WtnQg85wXwi6MV/0VtcAy8skD3YGpabvd8SOJgBjZ3GSQm
jxkuaOEqnmuZwlqOkyvEWmLQB5uizQ3YFsC1663iv8yi4mz2Vy0MwERNXpVOs/D+GGHyHezF67pv
9kZ0Z448SO2r+vRfemQ8mtDk5aVj1sypAn2QEiD7d11ZUSgt+1yZz1CVUHyX8uxQEj4ZPrxAHYI0
ScZ2O1fzMaWx3p2PAdEL/FLmXDmX1ZfRQ5pLRIjnU2H6WsnYeppD6qoFWiEYk9+qh55z0CRC6ciW
mUrqUvBmGHJnhOnDtua33XGb2wws3vNv6TWzrc3w+/6RqqMykqs3LAISFoeLXSVFpR7Xm/hd/GZc
N352WE/cIFCEdR/s3L04+sw1xMSvm+8l5VLNjD4xRnYZ0ZgOKQQBXI4LIK970MzimTcUKeljWb6W
t8rql8Wr3P4Rah+YWbD7HHbZD8q4PhdESoleTCDfX4Z4MJLUqX6ae2A1OQOTiyppw9BpsYfpb/NC
9K4T59X9EfwLum0OG8vr/Y9j7STtT6BkFagJChpuimnc64hoCdcVDP7Q1PegnbZSKd8Zj64F7XRJ
59YIEcTiEm4TqqKmW/SnJhLoHYVa5hoeGpF8bTimNC4Sy3pycGM6pMG5HjFI7tMWbDBOnZi3tL5D
2IbLiEhDxiq34q6X1vE8WTHsWRnnZMlSoAy3tvYJg+kEnEDQisuWTnEa0CvBhznQ2cUSvEW/D2Re
M4zDM1BdHam/elF9X2lo+AD2ZqEp8XHTtBO+w0MwvwU2ju/QboHvgx3m1K2NF4ygbvR2NcPJBLw+
f8hPedqSo6g8x2wurmdZ6fsZPPajwaNKz2i+TqqD9ocCxAJybMNm2usog/UerWnqllJylN2JZ1Z2
HOzsMqUO2jOWOq4hPRwAc9fheWuVmHQQeCecfraN3fKiNTRHe1NjBaKPp/eEnt2GcO2yH3pXpR50
s8Y5cwtk6JqVNTxDMYLqJka+PTH9cIh/P6fqKgFfGUDxQsCwrOnt5JSVvZsofa+WWFPGeLC2UpFq
94j/+66qryLtzt53BchuLOKxVfbJB05QleyaE1uRlW289Z5dHZ8AYw67CoIJh47rT4mhogiNE7NQ
c8dCggOANXWKc8g9tzEB7FGRpYCAgHZjRdoJBGtLVSG161ANKg2oKXMkvoJoh4VF0fOkw8YhLF6f
Jwv7svI5dlToJYF+YoGAJOvGPvq0QSDc3dfYodIdTtNtz3yZVNyETWR3Xdpz8l2abi4u723fRZXC
Dz5CIr8YJjicCkbELy3x1VFlmZhd17xVG0APC49BDOnCjXZEDJswoNPCKq3AahsfChxXug3Vs8bW
CbJAqpkd781hUOs5SrPetgp8mwwDcmvJL/X+rhaXWecXs/ZLTMdWyeDvPPanVvqJfF4C7s4eihXb
RveDkU4h9NR37etu7BG2M4w9OCZpa0GcjPReeXLfQKX5oXxfe6/U7H9yCdwctrhDf5u6J5Pq4d0S
1Hirz7fZ5hEfRH3pqgHfDtkcvEdsaCgo1eL3yTfrw8cpR1flJ4E2Cm/wv4uEjQG6N4A8PxTCNHqG
SqL+oty8iJ28UzB7AyAjLDaXa0uFMKsI523WgUhagunDxz28xQq2ufOvK9O5jwi5DWJ0D2sD90hO
sG5FBWJKZoK3U11VPs/JAiPyWCthdMf8LKXT/tYj2O/OxNd3+mpV4VEoB3sQkY9NYINjl67+Jfnd
hn1c1zH+iff4exnAeJ08H16jKOdAkYeOe8P5AwByD12oBDj1tkUD4d623UBqTmpflCgmTXLkzVOx
OctFiHNZs4Xad47nNQ/F26nqBNFk43oOdKtoXVQBodGzAWbV8k9edxzsR6Oepy9/G0Gk9dNeLTCj
IvXN9wJlBVwC0wYMvkjV9eyMr9zfK5BoPxXKUuhv3tw3L772V0kVLdxk2UdKM2IOO+eV4s2oxkGJ
sostQGZG1gEy0yjYfmmjRyoSFOrKQ+zjRjMazCjkFkCRoAEc913GXsbVC0T9QQ042vXFjy7GQX/0
4FCGFcCgkhLCpEE6WBek6UTvcHt3p4gs134uDa7msFtDGnXr5lcp7Bm9oQL7xPIb1iRbv44kuja5
oLOsmED/9M8KqofYkL6n3B3GC7WihCwt3zPRQOPfbpi2Awp1b/1po9lpm4sZu/nvFeGvJeOVWr+c
6GdM0QzBEkjmx1KjF7R0bOsC8++acs12ezHfxeJu7X+MM/TgXuJWsZINZ5mHuZ6Qn56lpVCHcicP
YpG/1YhRQoOLx/YNnhME2yIuCpGlkhUzEPnWbNGFf8cJKcYIkb3Mhcm2iTy2yQgacHKCjkI+vfJK
yKX8FuehIsdAdj4hpSw2g+Q66j8spqm69QXxHeq1kMcs6KmpnP4DVl7I5tkFUADs8PPJMdDGSr2H
a3KZaLZPaFZCooJR/UTJWL8z1Uh3aQ3EQteww24eFpz+iIzB0hdAoX4qH2QIhKwHvpVa+Us1wRZ4
LmEqSVxg/TfXd5eYi7brkLGxgvlWnE7nxJBvqQi+cvkBLIvbc3feipRgzJ8WTZr3DyARK9d9nCI5
/GWCu/S7/aputY6kcvQpAKsMCTiDP8KbC9MgzHPqisSuD7L1WRCwrtivUB339uxts9SJj8XvWUcl
rWgKko4/QC2GsymR/P4Bj9seFqGsjdXDPj7WcAuUzJsZXHRDbEBV+dB+Fc95dRUV8cUFaU56FUbJ
YXDRM1DEQViz0sPjrwtvbl61l75hu8ouQGIOCm36eWEabDWzaBy7EmUCCeVTzXWmJRfPuKB27Q8T
yT/Qom+SA1DT9stud4hgeor4CoU4ZR5zw71YBs1fPH7JFAZKALmhn4QE1V+fkQSyOq9p466IW+9H
JPpe4fTkDjKIndam5pobLmCTgVM3jpIhMXRU5WqgMYXQFn4M6hXhkK6MpjVnima7RaoW7AK2IoJ3
ZipXut35ViG1UF6tJdXO4XXJl/UYgpFynMlfBv2QhCha/ZZDw+iVLWjlcxPwlkxKqHJJxGRiT/TE
T0Jeng+DRdk55aQWgi49HO2o9oFLgCjQ2URN+OLusMQxc9XzMC5AA+wMB9o8j50torpQ+TwwKXB5
3+2SCRnXoSCNvFgejD6UvjTZtd2OwqlXg+78zRq0etwbAgo0iw6Q+widlbKXCo708dPrnJI/AcXn
QFmMnSRdZZ5+tkT4BRAaRxih5FuDBcKIEDHETdBKqcsP04hLw0Ed0XXDvYNjkiMFSyX/cZ9Z9WDS
m5dYGtCAi06WTHNWh1tZfDPwFp2R45EPmzRZkaCoCSq4hMr5q09WBdMtXgMpvHv39dCCXVVyGUcZ
OF2aDR+UVRcwnIsZcMr+mCZr3Ie/snRujz9i04yl8C/KaYpinH8/Cg/vhxlPFZJULjWdMW2mKP8P
qYxH1Qkp8zyAwRtD0UTQINQZ5BlswpfivLBuGHqIsnbjcqmP8Q/xqw4G9DbitiDTora67lzndoTg
MIc+USUDMyQ6nsZ3StrnVwMCWwBBeHz681J6ifca9ZT/nr0Sqq0acSPSHzZwdUrhMVFRDR8dbwyg
kL558xUP9pAEgslSkIgsohpvhF90o/tPjNF7Hd90ajVduw2ntby6RH4Jen9EGw3Vr/hgiDfjNq/7
QJrDe4TP7JDhW6CkrFgjTlkY+XKNrvuhsE+ZhpTNUVhQbKm9yVyDKvHkU5X2ccrsW6WSioJVqyyr
3GuVXYDrRhezx7x7pi0EWHC8a3T2komQ+wNK3zX4m9dmD0y4GUd/DEU32S5mGMmrfnkhrmZ6s8HE
2LKB/n5Mf0UFEuwcuWRBt0qYVKJDjAfehLRQPZFKutiY2ir3No7Nb+4WeMaStkIgmvzC4HnBjucN
fJ12CnsQ2LaOpmMtjX71B/Wpe1xXeeWW6iPBEP4U9RlL7fi2QL6YiW8Degdtf/4rHb9ezRr34iXX
oWLpATteN6SIV8QZbUQ9WSnetO+L7JC6CX/imUDBkqh32Frm/HTgMW89AsXt4geZGKGW8PGajpb6
KRwoa0ApSqTvwHk0NgzG6BCAvq/zwz/rp6LJZ9lQ8vDQKhSSG5p8w+0JmAnVjoqk6twiO4F0ef8r
i38sVgbYz1fR6oPDSH4D2m+H+qzKmuvyDydLnQrxgj0jCL0SdEAl0gjyWPofV/duF2OoBqH2S+4B
HXMpc3IIQnfiGeFoPakYEC5gl4OV/bkeYNiNZBSJFjege2QHXxcD1+SV4IMig9+0RSgvLX+tho6o
E1yhV2QanSGVonbnuNhHqNk+JRpEoVWI3lnF7/LpGaE2zx7Krvv6l/GyCujQABfrx307NV8nWuLq
kuxE52pHeQtY3vu9CLampzGtAwRpA4BD6vIPx0/pR+VajCYiqd1ghebZlM96fucws8Zh6VrR7MTW
6EA3AcqaZp8pECR2SicMFSYbun+bJ2CRpW+P27KtLvZKhY9V2syCd3aSiZbswXTYyPBkoWL1IsSk
o83HMBh4uQ3zqj+JLupZI3pK+2U39YwBnNiESY0CHXUfm/6P8aA/+qqeq6OlKYuDPXhWpo56L/7q
wK0Qmuw6Q9EkVSPBYal94LnMypQJP4v5P/1BAzgllNgBMlYZ5KbuQyRLK+vSZ6LxySgiAd7NPjxt
jp2IWJu2dES929V+RIZcqneJijZCz+mUeQmJ7Ag7Za+CESIJjfMrH/ceXvHeqm978HUwWAy8hHY9
e5na6BRu5GpP36pl11vJKx0Wf5mJ0Tg3KD88Ajh2B11hckR4dY7V0si3ILFCwa1M6wcnmmLaUKrs
Op+f1zN/fdfqTpZekxBw2kpvjXhq3qHo6r0tgaPcu440fVGLQt7DGMJqt9vFYo/crzSN6bfVbOrc
+6dTGdY6c6WiVcIsynxzhlaZUveNDBfFCdhFm9GFuBCt5ADQFev20EU20AkxF1fNY2ln9OXnVYBl
fcvLaj6NDux8HzBUVqb0JNLquD/nm8QPUJHrP/cSdkOnj264Yfx4itcwmQrYMIGBzwYSjXfXRRsZ
apI0bft4BIxfSpU5iSZSOy+BDVCR1iD6dooo0Y5FJf1dDXn4swPKw87kWDtElmxRvJHlaelumzF6
xBd2jsExTdHVfSoCc++ygqlmnEdCxKSuEAmFrpRMCP5pYGYu0hCBh5I/MBMSWKqu3wBJsxbHRbTQ
PVyT4LytoFLPZEMVSDrp5k2mGTlcNrK1DW/CHPofdKhPEcDozmU6CONMTXIsCZDfgmDqVyZJxsxx
VcwfEi7uZ2l6+2GTEis4BTFgNZvYv0Wxmo20HD3VawC0PXbAYunA5UpvLFg4HohQswD/Fiu3q6PP
XcY08NGjgXg+LKzdaA8dZDi+RwsYPiZicOKCJe+HVeU5UfXLwAqqqgcCe1M93qyro6Jnq18f+Ehl
tXestQOu9HrCGOs1yX+IYoleSiXfnpWhoCoOQCaUBdgRtdGPGuVyyud98JOQVPBjvy+BDOaVkFAK
D73PxsftSsybGusmlX/RutW9MNQlCo7EiLkJn3Mil8TC9vM/Tfqdovf3gjKYutypz+BZzKQkeS+2
H/5eHeaw92fRMjR9I5rBBQIjne3nWghDgLaOloIrn6cMAbCH95glXaMOchlnnzJuCe5LuJcw9HXw
77yh+aqeQYYVDbLs/Z6dhdmZvnBlkjKtL7DJx6zKK2ywML0Lmdgz1SU+/w3OHrezwf/DeBIsrdjt
4fVKov4gBND0RmZYhMhSLRqu6BQapURqwbdmTRl3hwUedyfavtgAvh0VEE6C/k6+6Rx1RuItms2q
D00bO7+jkNDeV1OhOY1rGqh18/mx9c7WEr/INFCAy7W4j4Fh9IaW8MbkQQXxZ8eBq776lwWnNVmO
n8KAOffzvkKt64eioHkQEURoabJD17Nyl0+Mhn20kZCNPt6/be+HAJRcnxE2vNUTmqdtMjAwHuP/
e2QORkz8tFDg3cT4hIkwngcn1i9VJ00Rp5QdxN9Agd4QjRq2t5QAdhT6axnowdObhk6JB1E6YakX
4+w8aSVPMUsfgba6GfFMLCXV7g2x7e5kLdPXBKSPIeuBqYj9EOmQr2g5TfA64LAFLNZ5Za3npXtX
xMOIAhsiT9h9JjI+EXZbjDWgqZEcuI0hQ4WrPfrSV9rnS8sQ9qBlNv76FdOBQDJHtOZDPbCU8t0O
YZDvCGbcOXYtO4vSCD8p62HDdg6B4Nlb8JcVKU58dSUu5P9vFOdkxJsTXXbdh95jfjwoyGSE8XBn
oFXaWBiTe5XvfG/U4lIqvijnwzQLzb0LmKnOhlwnE73aEWQQh3NRxTzzqBB+XC0M9poVADAhfxMv
vS7SqHziJGOfRXtptA2efeRr2y0nFwAXjAJGbPvIq0Em9k2aExNkkGoVZxiPyB05vclL7tmiP7E3
5Xv+W+eql1+10vVxyCxQ9imOI/snRMfgK8PmDac5k+VL5mRhbfzrlhspXY52phdwblp1RgbSsa9a
Ujg0LS3fRauezv4i6/6wLQ9g2EqENiqk08PudZiaQpotZLviYLuP1Bop4/R/AWAs7NfGkMzVfB9m
oVZNvZv2YueEC3vcrIVMc5qlWRyciQT6C/sm+fodPkKNxEM8X7OUuKZrX7/QYsK6OVX0qA4npexo
avYzS0zE3la9ZUPvi4yEmeEuCWk8o5upt/OoNJaAyfLnNOlv0ZuJr2cVROoKGEAgL964UXXyYz9Z
NmfRoM9+Lwf/K8Y0QnthP1tknb2Z+E+TXp3TBqDpckh1lSc/GSf+gNlwa1/NpVLX5rUJhlbGSMZf
1rOM6Pts42wDNXPt/b6NRWaDmvFZfGUAhqdxSnRA5hS1AXDVnjG9QFgmCBMsSL/wYSdBh0Dt4XZt
F0gchP7g+EJ7/KIw6Oyor7hGC3+zs9tPrfmhm87/LyTiHVSOIKaE/g+I52dDFkZw5Tf3+yFi1pxE
1ywwQImW8BoWtxBGpQ1no2KRE2wNbiwBGEGIBhHpMkZUOkBhRaNAjbgybeK2Yxz0CBZCOEb699Dh
MMiRMMN7S1fxRe6jPyHRat4n0K7vi8HPEn0v3VPlzeQJF2KFDn1cS0+IZ7OCxMCglMXBabCgNhHw
3cE8cwJ7cRKtKj/yLyrhbmNjqQx9KchxMHz9vbGnI5D75pNlnwlOuctv0rt66nk8NBbJ1UBGs/QG
I5551oLI6u2Ybd+1e5u1odxjpLx2gXJMl1tcWZx7MbzpA9qMRvxHBP/D/+gWaSz1F7tYTzJuH2sd
mNRHOGMCv4TxNBm5SPHnlnnBJzxbjwzNY22z8XlFaR1AFaqG88r4YagDVQsp/uRTXmpzcnxBN1SC
7593EBGS9iWrpO1Yyjb8sdYv4E0fARi83nwncrUbwEDS1HLu7o6TxMsCiPJzevPKHIrQjChZbJ1S
cq4HL1FCOk/8j9QfX4sPTSPRQ2C87eA2w3v0pEjgiUgPUSKS1zI9y0i1oMfbTcWo1GViP0YhIZb7
3GsV6Ui54NMPyb6bCz4nZuxZauR0Q+InGKPGEDDK9xSaMXJISa1TCkYvkVf8OKsCPn2YmkxUWLP2
hEHHkNXYwUHgRwvH5QVGx4m0KiNx1FmIllQrHivNuwIAaS7nhCCYNvQNbGa0EnEe+Q9hrxDQto7Z
QbDghIMplmZJwjnZ1WuCSvBcyD7+SjqkOZSTQpytQXEdUE5r+jQnSLgca375euDeHlQJR5QQfjTq
wCkprPkf8dEm7EYk+Y4jD2uxBdltIDxO5CIwpVqZ5dnNljVpAtMQFvvUM957csswVQzpTxN1md0T
o3gfwG6kIYWXmxIjIotI2dP5QoFL3Q/2oCeReu1mElPZA8n2DN0nPmIT+99+4ag/C7bYc1E7MmWU
JioYa+cO4mlN9dcvCiOynu9EobsPnjhAKY2Owela/sboLMNhLRrNZ8jlB3ktz4LM3jybO1f+42vb
ibdLxhI8fxBLAch4ZTscikUQtz+wR/U4kL5R3moyTijfhvvySJCCHEkvx+BEaIJVL+XfJYRzNn6u
j9WvCqXHU2Rhz9GyyvZl3wpsoHnt8WX9wxaDngv0qPyLUJ/Cmko/ye6R2RQV96DEmqzYelXTQf3U
lRax541sEsJolJRWUeg/BPxF8Bn2jC6pshdizHs90ctOOru8gvLXxldUxQ7hUGswMzscj3SzH308
wqfporO1BI4E1AAvccd883XIZ0ZWmqCMBDcC2uSZi9JdhNIgUT9F0PhyAk0j39YfF0nkuZkr7oMu
Zm2TJosQLb7//2QV9UZJbTlENPxuGVLJGoSKxScMRooNua/2a5QpuDN6qft/bfQK8uglOz2M4vbF
RFQQvKTwSF6PapUBmnRKuDHAD1FMqfKupTEOctH95FID2tG+NM7//I/m+VONEdYTjkAQlawl6A3t
StMg9k+3bwQJ9E/QcmUiix/VSpqQvrdlN/a/MAfpodncQGHRtXe9wI0HHQgwuSV9cb8ngk1M/4SV
DcgUiC2H/2pxFTcZ9Gzj2Sr5OuBAnBhxO6igweUPxtpP85RetYMIlSqskUe/5DDrDvd7IGRNiMgF
kG+3MkdQMUaC9rE5lzdBQKyUXErTnCg4nxhMUWiLC0pNV/9qaHrMYXTbjoypla0PE30cEh7XcJAN
wLV/SOFvR1f1VU/h9i0b7c8rJ1F/l+4tk2RX5VMSiz6FX8rJZZFUG33atOXJsJrkXtXrm6naNdpA
bSqxdw5f1vmwBOD87f5zGZ1npZesvjcqN4BDGhyrNIl15gbMOXxhPmi45umHiQrjygNnunEj5iWF
DkYvr8rUbxbAk0dJb55S7gxhQV1LEjcTfy9zJFrjui//ut9GbClLUGyAszPXaRS+l2AUeYRRgu7t
WWnWT50IrLG9RFdlFZNP7HweBuNJuFMSGpTqnkLqHHEvGn5LcHFLwhhGgF342NhPLdPpJiXjWGfz
+3YcQbVqd9me3K3f+uCAXt1NmGrl/QZIam/8R2TTEO2B+lNska3Vjqosw7jGB1d7t0c8RO+7Zq05
yXOEyPI8bV7dukbOLzrfLOathLw4nnPjlP5ZWmupo7RfhihkyDGbk8NNuyCUEZjZbNDy8mywRtj2
ixjaT5LUvieiNobBzRIFiObYWB9rw9HzcysqzdTO+HjTVn6u23mh0oyzF31kM1a3ZHek6IjLgdp0
6PStCmbtlgdKaNSo6QEZH0McNTkFe/+qhuFdHpv543312grBPjEoSujyTndae3iHMbDJvy+Arp+4
Af2rvxiMvUnUBWgOQQwamVOBtL2+CydpWITUIf+FtmCBBKA3ToIky7EXzbv+HzUNyu17S3GNdlAk
2B7qzIYTFRRAg6uQ/i8BuEdEH0gwjtSO/Ljjmx8r4zF/D3t9kas+TL5wWlyiWRG9jUDGRP6/083V
In/BbbR8aXJyn1w9nomJV2SONK/TXYxAnWx3MAc72BNdkWDSCaZyFmW/btYh/4AqVY9CnOmYUujI
ns3yBwUUxOh4YzNVI2PWOGhpmJgAepDtpC+8WJmLlvUAyTpkUId9goY34u5ZQYlPAGWBC+FLrI4V
6mpSjXU9monxx9ZUk1dJtCmV5SViYYTs9VEs9RFMCWtcBGaTD0FfsCJCBHj1MclS+7Fsg3tpIsZO
XULluK806dhGF/1OjO6RAKxy4bU6uMUdJPcB5n6efzQBztscMSBuMMdjjAmHNbKwP7D+IueFMDU+
OCWnnNEg1Z9xisTMcmHjX290JXglOTzZDKJFE3LLNdg9kImQ+rzls4FKPOM8iLQfJU6d/FpzVrbs
IRH6bpcMlB/zFcrc07blhHUEW8snG8KgJqiowSn5R31JNXOANlMNsxKAkrk62iPKc86V2zUcJqE1
ImACvpnPl44BrBmLpddx7Ur98oHGTcFodQrCSG73rcD7XNM5xPEKqkDsDdiUo35KHriKByuddAdu
M79F6XwDEBtOg8tyaDNQ+bAplEIG3+sfafh8Gdr2wZbXri+L/5/hhiZ+e4jgW/IyG8hWATnbjqKG
Dz9iai++JjZIfEEE6nRWpjbymecRWwqULDvi34s/FDXV0jMi2aVVoU33oYY8XIHZxC0MsrT5UPuY
sZkS7yKibIRram8D5OWRBLC/E119fSPYFK+0l0DzrKWiNGWQRjb9mwJ1WoyJ2ygHykjrH7J3olJb
Pwmkkyisd3rakqQCDhwD/DNokPTA+FvLvPs7D0fQq6UegUf03bLtV7xKavSF1WB7PeKRhHj5tw7X
BGhK2JW/FAgZUx4CpaaTUt5DauggQTUcjhEf7hDz9w5nA+pnNH4+wVCO6G2nuKo7wwNJVDlh7zs8
kxXq4MINMfbXVIQ/xOPLFWbOrT2dXaCPh37yvZUsNl91c71sW57vzYdFaOPd3b4JB5abXtlqVsfL
85ILZHMjCjotEKHPzoQCWLE1A3gTUAaeX70fUAedFB4Ja+1Fc/VQy4ldRGGd5ts0tMNUtJ8SMYuE
Lim+VwyS8YT3rR62YV0oAllJZ4i07Mjc7AnbBk1u3w2oMJlnz9hHq/WoXDx/yEWxOgCuFtAWTV+8
NxGY9xJQe1q7CC3j/F8kNRQ4pjFby5ilLqVrz6u2+aBRA4IC3cagzr7s71pCud1B1BmDEmV8rFXs
XrNSP8xOC5liOsru44qqDs6kOj64FK5ruTsidv/WSan5cNW008c8ch56VU8oD1QdnGC70zYqAvtN
Zal75dxo1EmvllQnv/qI9lezsMOYEa5DcM5gpEJWlVjxiPmeHoQi4+QMk+Ef4S+tarwVrXgiNpjc
7LHwMSI3LNPZ2Fmh8lmum8kjsQtLF0XmJ0OcpvybSKvRRlOXS/VKy19ukMyPXzhwcrf01YRytfmJ
JNbkAx1310i9fR4G6i6vpK2WTGIUMkwd8W/X0GAZKD5iEPQU6/bsNDnbQo+D51aaOohA3+pM3bae
GLeSBg/4iL3E+aod5iNyLRrjIx76jgx4zq0ZwetSnHZAhQOOxxvvXN8j8nURuh9+QzMcLP/K263d
83i7lzNzyIg7XSyjXfe/Vj8qR4nd+3qmAyaZcH22JJOEw8L7oz6B/cN9tD/ksNwgWH26GRwkeUQk
2zJ7JOr49+ufTPuailkBY+HClQc1PtDMRd936JM/sQnFVK5RqAMUokIgCUdpheIC73lxV7NqSYEr
Ir8zkVJVI2mqSXs9h9TO5dlE8TgUwjwI3dSj/TiuzsY8b+CS0FdtbjQEjZtux1KCaxBAxtMcX/Zr
lJ5qKQBK7URsOoTs8eUyr4Q+5ahhLPF0at9w2dl1bfAfBzeGgzx6FMat84/5g7tPgvLuIekzNZz4
WiUG9YDyCTBYlYImOtRMsLdJgT7SIGbUBOSDrZ2XSScZo5N3Jzfq/g2uOi8NHS1O9QgY6wrIZXoR
IXQh6TCGNQF1silOVU8kQK5vd/DpMepm6NKMaaGuIl6qbz5LaCF5Qh/JKWx6sHVaLuCYXVcqXSP2
9KXSgSMu/+k9gPXjIv9R9oU8p/Z5OhCZ2sxlLOYcueBQXW17mSfMECAe5Xl/x7CO/AMJw2liQfhI
B/7azbLb/fK7i5SYZ2eIQ9jpHK0oA96/5fzoMuvZnOQDgFAzd4EPdVjdMkvD/LiblX9dr8mNboPw
JD0mtjwwN5Oja/v2/BbgNIYEXkliVstB/kUJ8dftZViyy3JzhyiOpJmDWl7Qyzq8vjIV5qpAYNEm
OFR+nb6ckfmEqN0Og6jLrQCbOD2aGHah6VuYOvuq9CGmOHXM5rzoY0Tm7xxaQkYTBfRyoKNuvZld
oJZ5xVpXiWRBNHGP43OSl3Vul6iVREqn6bRxLw4ke3WMPAvRllioPhMgltiLcJtJTCwCIoy9n9PA
h2VKDlPDKGrd/IhRUscB4Isuz3W9xs1xDKRYnwR0M18qcPjQcDI4ZSHvVQ7TfKCwjj1lVptdX0rp
QLZAaivrISWKxIE7RSoVSPO2FhepgUfH42XRfjCwQ6UV0G+0NNlIAD3T0pz2vPsYjzSNW+orlMdD
PE8CKAWl+DTuRr740g7i7XaJPriTMRul6V9bbD3G7bcE0qRHFKidJ8wgkd6FtrO+9WXQPGas1GSO
JEc14+uPGA9oLr5PqmlmBPNBOAPXZ/loin7NMX43qSKQxINRHzV6oDhgdGzjLup2TcXOSNW++Ljf
A5hnJugOdsy6VvjUnFKGqB2Hk+zgC5aDHY/YDVS9eYps857pIbHcPRWPS/GHtwJFeRgOqrDQXPma
SI/jxiT6TF7PNFf4nvIkU81r8KN6n7l9TRhQRCoU3Bq0uadxlRid/xsogXD6WbGv1RVo91Q+TlNI
KaZFMpDYK8cqvo6PuQmciR11AcR5Gm/TiJ6t3cKNsvjypX6qlZhRhsUm5POZOrguOcIx/n5nW2eb
RK97LMjpFhc96KckayQvLJVSIpxSd0Ar0Yl2PhdZM8B8tYSM6Boci8dlmk5s0ax1EdROTu3rR1fh
MmTQWFpPicz/6dl03t0MbGf+fM6k2tRubMb2T4gl6nfOnxUoN9Lo7bxlV9cyhyX+2GJG2EsObYu2
1Y4jIlBBFUdRqjwsGq7CiwsZqNifdANLhO6Gk2xNcD06DWGPlq093iVYAKB40VlkCFbIHw3UGsp/
wsWVp8zL3N7I9tmIP5snEdhJ8UFvLXXsOxip1vC8Kt2PUT+H4IMoSb+Raql8rcGmqUASlbBZzs6u
WW0AYC2UHdDNIcO3HeyAYYy13iwsE1uMtKxL1yN1LaPsWW2iAsKwV/lbvF8HRBSy3A3ft6MIosZJ
rp0kBQQ8WrzoWt5CI2rSz7A8N3n1iNIQlZINSby/fkBcd70WlgSQ26wlYoR0hBshFwTK8m8NUI02
JnXp6/g4b5bhL/DwStWmEvE1BuhNEeOTtr6+7SzqMf1iuFyyrGoCgaoLyYRrX0Q2xBTXttbtDGQ/
OuCxw01H08XsmXKHkK0ZbdsAFFaWB557NFDZs68uTT2kLzYcUZsddNci8HDn+yFMFBjpN/yfhndt
fFxXAJqlg/eELOMvG/l2Ekiq4mAcW0TdStKuHp4qWlkOttjMi1OGOE4SnrJd4HQZQoml4lIlB4QU
2Bi6IpW4Cg9wLkBHfP/EJBboOqqRCy7R1zF7sE9TYRHNjZaTyLIa3XamCwPm/3XlIKZcNCMAucft
a0EEXjSGt39WwNeTSXK0id7Fy8McTbY9ifDWTtuSRXdre6MtSiWCjRDKRcT/5jY+G4lbFiU6UGjw
4dC9pw4O9I0tqKCHzm/3KW9CE0vOKkN6sE+mfNwbkUMMkXm25CLut5RBelRTQLKJEG0jxidPse7y
s62Y2oTbVQzvD0gVa5T4NOm5XK4OSHX2qIbZ+oy/G8VOmiuhDmV2ua9MiR8xP7Kqk/y/W1BJVe+Q
GkyKXaK50/datkU7m9OK7trrbpgTkF9mbLUxvQqHkB2zrfEi3OkkVWX6swr4rDkiUX3C55fl334l
+B17TlsksE9MufJMXm+XnqmE979iXtvf536H9Nk1sFbuPfbs6LnJoysIxQbpKBv3VEfgPkKn1u2O
16fzxtSLet14lhOLgTCZESs5UpN59DaqZ5EtJMRCR3dOoxI+dIdWsXVZ6ZMvXdZx/h8JHgT2uCyw
SVNjT8cuMVSJKcdCSJZs+8zzVFrObUbBQA+CXd8jbGfG6/HKyqFl6QPqqQZYy0ttZRGefohuW6/K
HEuQUfHuZoLgMoCfVV2oaOl+6QULix+OGjCgqR859NwvA15w30HEEeMyWDyl4LTmLUsRYPKupECh
8dMVRY8l7NWSNyDH53d0QllhwsQ9xlGT99M7HZ+12E6FTu9xVm59DlHocQWzD15FKPSipO4JMY2a
vEZ+nLJIS5nvwllUJb0aehkNFF1SKsJDxE4RhVf1HLxmGBQfT2woFVK1aau2+qhUKs37Q21jh/q2
Zi97wCrTPoE5ntCkjpkL/NaSd5D/modecfy+NJX7MJDK3CLw+NYBDt0qi6UmnoUEYJwaNW1lumM6
OrQKs7d4VabXZFxa7ksMAtozeyL4UpdHfm8Swjj83+SUzOzRRSOffPqfvXWW/1I6TTimWbt/n4/t
XkT/YGL8/uq7A2f7B7Yr4lWnamXoIj9sqwXxqQ8HMcz3Em2uuNj5KJfBmKSqBIMcIC0QyyM4O9Y1
ErvmMqz6yIHHvA3VugTKF6jMQ9cTSFpSHOm9JBXSW2ZmD2mrttyZLEC2GCLTdGDldSF2jmoGQd75
0Ssb3uD8WudONC/3YH+L9ia0sBZlF4WGbsisI0Fpjy4beSsfVF8Rd2YbNHIffLv7FLI5iFTWtPzi
OBeBbIdumSBCNjW0X/nCxVkpfRNYcoBHumu7Hl6vZe7C4rLK6qbKhadoJZ2vU+6xsUqP9TrWDBhk
JvjU795hmvRDBovgzfzk2+CcoooZ0QdewmxnmEbQSZuNk1isTu8GroFebz/lLhbwqN0O7924YZ3i
aJh5eP8lWH8Xx4pcs4ojz2bQrJ3wSWMvHC81doHcJsul5p0Afd1btf9NVaVWzDbGkjyb/BBIlVNL
xr7CNn/Fy4bX7n9OIBtCKxqcvIAH9STn/4T/nnWlz+Mr1h7MZY21uNHiex5Jxa2UOV5VmoMGyVoN
Ko4m6ehcoEq/qQnj5eGUO7F2N0xWw0MIJ1lDO00aHKo23t4JAQikclEaf+wEEkYOd3ZBzkijg1QJ
WCp+hUEySLFcaMiLDewIKoK7BxWHR89DQksHzo3BMPejePDmtVK/fjRkPIUzCFxrmkslt165kZ7b
mGyNw4xsoyMMdaDbrMTykwugr80M8zzlfYa4W82IcWxYShdfZ6sq/Ef5WhrhNIGm2Gm5b+WYHyoJ
RjDkOb3bkGkqI/dYroidNAlJu25W6FN0qqZ05NVI6uYYD6Mm81RC1sI3JBEjJL42s9sMGXWuqbz2
5kj0e6dHnzUOmsujILorcZppWvMEzohziz2XB4Tic7jDQncUzAJiQ1DT5QLqtsYDA/eEsXO+M/H6
8/EU24sQDVDnApt2fUvg/8Jm4GCLXRlmPqDzy1GS1wzuPSdES6L3YVQcl35xLs9R0qn7UxiLUk6S
THmE46nmYkYkmwIVfHSzTPCJe29JLwKJLGFZQxW9GaB3Suka4fAKJecAuV0JuMDeEGs8nhHh1cCY
mNn6pyF7BS7vwUf9bvxhCgs4+VvuxHJCsg7x1UHfLnpDofK15HWpOpYJ2B7GDS3+YCGmkfGLbmcX
vm7QBgewFgGAxFg2tg9apwDvOlhKs34ExpkErBhtviUmcL0ctM6EDD1Wzej4xeh2M2xm3A+wEevA
Exo85ULayP8lq4rx74Z2oF/K6EF2m+eXlC6uKw8IoNz2PoHaIhYtp+9AE3nOH1yToF9uhFwUqWbv
ht6o8u7RrTPFhRXqJXCSJ9Ar/VoHbg74KQjz8rc9M/8ay6gbRoGcB2sLZ1ZOxwtSEXHBVB9UaWTN
OmghOz2+fqA8aBQSuxKNym3bwUqfnRTdXUpcBgIgGuZ3yiISy4FYegIf5Q/7VUe1xZ4/EESJCHFQ
FpZ4HWqR4H0wXFjaYry7TbKmVQDuKLAIW0nja7b04juRkUIKf5W5an/ch9jcdYF+zzK3Q9+fXwuk
Pg9+4OjvzDuL6qp/TSeEhVfKSOskuIdX23XZg3jaRY80oZdJLsAnwv8y8PnluvD9087Zxk7tZw2a
9Vqt5YDv5FWXa30pM721F7aasma+1TAYR0v8euskIATKGodrbUT+iUiggfDxm7pEZ0Uoloi99MTL
0ytgwsmxCvkOMUUscH6yaMZgJ4pUJmXMBFgC47RRB61jFHJ1Q5WPo4tFIb0OYPeCkr/oLJA9fV4G
a5c/au1Lk5EkjxL/Yutc7KBWg6mlNU6FAQ/OOq43zrKUTBg+DhZWmgvyXIIyG6G63ABZRHrMDkUS
pJomxw3Wc4k0/wwKS8CbeU9wHM/uHHkgdu0HPDCMihdulavs/5JOiGagsp54n4e2yr6IpuvuhbfR
gbrwfgrFlq12J9FZUCLMYr7VN1Cv4GNM1GXcnf63Jqb9pIvsNxXNgec5AcWgoy3vz4OWKxXaHlTT
ynyzip8yDLGcqHuc/rexaT169y3vJSAN86RqBFree2CKnF3HP5hbfL0LwI3s8qfwt0U9WCTss8z4
g4ZXwBjUrRhBKqegrfeYnwrx4cKLhOy0YLsoVH3C1y6NNYXb1iCfMv94J9gWfKBT3V2l8H+LgZ6d
dBKNUcyqT1lCxQ9VMUcG1IX4kZQYvLTQ5w5HCciV5myWYEfU3hPFrial6lUXyrR72S/w/iZCyBSt
2JsgJd7MvGRDum3hnPXt8hDid7JOG7Ri0Rp6hd93FK/6uQ9JopvbZI1U2MpxgLiQ4eB/xvf7LsRH
4PfflVMPlZDiu+7rQ6SdNDd+lV0Ukn8y0x0/3CGEbGLE+P3lArMmEwVQc3vzzxoSlGLY+X9HyFvH
O7aEpa5wW5Ct2iAtXXLEhM9b3ohAEZqXNbPEzPQfYrKLIRDdwBOwgAdh0eIhRLxbHhAbSMKkqRhD
DoAPPG/TvSrR5GEwwp3zmUJRMIWHhfYbJHvHd1B+q3VAeQHNsrImoOoiIyhS2QhQ6TOfzqLm5Z6D
yI+iKgRW9izNFTRSJp4e+hCIA9Auv0efilnMIUc8MDPKQ55WV43Gh8oIDnduLUDEwzMbjE2H51iM
cUo4Zmk9DLxBr8zfrI27x1ZViJN4Y5su7On24kd37TzK2n1OvV4J8Rf9/p6c6nWI99BrKadkUx7f
T/nIQwEZ83NwI8XdLB3DN2dz/c5I109wjSBqW/rTwP8P3zvqEIF5rUEUcJ6VOSbYIw50ngSM2zpE
yrnAGYK4bU/1GmgbkL7B93ovfFtfEX9MRZi4N6DGMazKNxOAbVHny03pLmrz/Fd1D9ReJTAB9Pwk
fI2Ok5Px25f0tmMxK3xMxeVDq6Vqf/zZmADbWh84FmrMpx2a1IC7XRB4ho57Ss04rRw96Kex6Jky
FKa++dxVNKhlhWKHoUpJwJ4HeJRyZYt9skcbSfi5sQSr7PTAYix0xnW3Plr7veGgo/LxiW+ZPOkr
DpqTQDfJT9yzE/vX2WsBGQVRyeiLLfE/xLqhU+avShg2eKWxHaFto3VJNuRTfW6kym9mjwfP7JxR
vf/QeOjVzxlZRLfupUACTbutpi8+jdefjIO78V5bnnv//itzn4PdrzlP2BbgWyfGaZAdMnkHBcTn
NovuQ1x1lIX01gtfKTDLYk2LokEEW2MaHBwGgKwyUejhrjeY2M2PBGCbGRZLgTRKnpul75OSZkYF
yZXV7q9ZikGtTw0lDli5fc9T2myBgAXBr7YunQVEUgMRvynMiFTDX/5Qp5KcQ067LnoSWfgYt2Q4
AEdN9I4XmRd83Lw0bkOS93CKA0tYNBtn/Y+XmHFJot1baeVk+sm514hxHofyLwru40e7toSJOtNS
MXaUFRLCPnjq7rx7w5kPkRvP4gERU9WhZRd1LiCnJL9Tp5+ovlzn1ahjok2vpb0k6ja98Fq2wnJf
/8zPjWNBSZSFi+JEl0gtn8Dnpc7B4s7nCqM/dhki39dWs5VrPJqwSwPLuXulmWpct+4kebnofHdN
f7sLA41fgCviR7lvXWtoTP4aHEe+Zy7KtbCjG3Ks4kwsKGdVhzS8hs6GjUIzBuVAxy5Y5hKdLJb6
F5Tx8HE1Gt8GO1PAm+1VM+KWiuJxHKi4h1vbxi7Y0Z69uz2hzfWfKAUFzkPK9k/kdoeg2YWYkEpx
6HCzvRXzUC4QUiyg+pkcAWdiIsX9YuL4b5w9Tx7KIqPC/KvzRB4f0ga/u3FDEgreIMLCXoubnIsY
0xT+9t9YmaPG5Ke5H4Mxe1Fkft+Etz71cd9HKFfLUYab890psq2gcqVBNuMWU2/PDuxq2jn2lXsd
ykNrUcMrT0wsBozIa/eHDvZSvoT8eYfCcTY9EKAnVfHxNDDoWIVwYGkj1E5dMlRQjhtnFs+LbKZO
qWbBlmoDmf5vgFMqGsHRb92ub0a0zqw6EC1YTPTSR8nWeLoSK/lNU045+uvsCI6/IzrlQCL/fttE
+wSUP8odTn21nBe4cBPJnE2F7ObdEAmFBcn7KSRC35zM60huXAtoai9qGFlxPJkG9ghwhj8+7hsC
llqbQSC8jPSDBSdVyRxPzH0MZ7ehgDvLzVNjfU158pda+yPyKutkBMMp45sWDZ7D2QqJzM9GTK7/
PZrls20ZH6J9kQsxW8+F8K2Knfz29CZE/6Ep+bOoqcXCj4mGYWV6j3kpoP7hJBqF7PKh8riwCwPA
wIC0A8ZZjIHDks2K1UB4c4aCexF4PwavWcMN8rbzmczy+aD4kwU1rH+osxokObXmdQfSAGoo4Ee/
kDkBgr03H55J2hxtEDRKWnbw/nwCpcA38HadKQ4nZxMaK5GB08YWrKWEBJxDdqGQtToVQNAcBlgK
DxgR3+CsScfeZXsyIP5mQS+wQMSXhOO5Zd4gH/xBe4+WTnf0NMnUHo+gaNeR3o7ZFF3hgUEPZ5kc
WkOnIh5ADZNt/9esT/wdW/UxlHdakKk+bc5OiDlSJnM7yQmPK2cmZOes9NTgS8S8tMBxeTfuqBvk
y078Hswhxc9r7WyRGwuIutgetHsz5ynOIRkXA7w3kXHtvELZN2rBGBWxPc7FJOZpjDBPit+LGTMK
CHIE9jazeAYaGbwt1NpHoXMNzPrB0R5ISKjaKxq4E1ak4jsu6lyUi3/CDarGVmNRJGf1eG6zs6Yi
1qK3jzLk8LKAL7A3dEEQbuURcqxnXEPzoUtDV6uJA87aYwwW0IJi4Ks4SV/uy4ytnJ0YqJF6ATNd
JGh8idpCb+CAaTcyEt/WZO+hcpuTANMmrRxE1I7Or/4tcUnmjcMKUo3mjtytlRLOZUh0e5ESfFnD
WgyKsHZj/xy4FjprVUH5T47YfyV/wDgOKbU4w48lPKWlm3HQ9Y9Hf+o0Ft6PSt3eNuhxgUSLpNvi
su0v1szaaQXFnqeXt1SrXqw7+yPqEtCpJaoYlUeWvNrinXNiH8ZD98ys39wFSK3/OZd4I6cpBTKV
IJLkeoFJlqdaZ4VwI5EBdd7ZdkBJ3tvxQ56Ecpbp0YZnSVR60oR8gb2FNmQ5T4jGPelWbOC3Ghb7
bYfsQr+bHSIHRjOCcgADIfoZOdlXgelgkE10uUX/upyurSbfHQ36D54lZTOC04niVIwFhdlmgStp
MO8ORO75D8dzrtI7YP5/G7NYvlI/RdmZh2ypUWCMqXzjoC6ci1ff7QuTanmCrcwjPivUmRkhc6k7
BFuO4VwAYc5iY6cmIrBKhnzlA4q5efL2g+/PyJTDpqNmRFASiQwlcQP3PAxFvD1JhWUh3MlAajCV
nnb5HzB1g/9Xq+iaVXm177JP1rNLTnaxNFR3bE4zom8BIUoUEVjWJnr9sob9mv9cJHKbsjfEPY7H
fILonNvItr1u2iHERclvsiwwvXpOiPWOheC8VEtvO2gKqNfWuBs8kS2YNJA0kWPEXZ0zp+xKbJat
6ktkpEPR/mHNVrY9c5P5GDTFV9Jqej65v1Z+eFddnTvcJosdAUfTrGZKXPL26F840gEfj1GibPWU
6LMrFMkEZ5B56+LMzECPYE6K1VXitdzTN4H7ie05EXvQIkq++IEwdBu1Q/Vu2VrmzlqLMDRIFjop
ImX/y5mr7kHMnSG1TsaTMpbkgeURbYSKGr1cc52OB9UaS8ZbuNwDi3hTULBo74mUFilUMHCYZxyi
ncfUyKhX/keZbNUx7HmhTgWtz3ab9mUMl2+rNFMpdsno8sYUDks/Ns4E5h9A8gtyQdX89Q6rZF87
oBUes0yIE9ECSyKBaFiUpjE9UnnGItku5hDwxKM/CUaUoUbfuKBLueGIT3upu1s4Nis5SxHqvzih
gngz5NvoRX3fjXcW2pY2dZFGz4GlCtJhYuO7g3OZ7KtpqaWrSre7QbDveVqIuHVmCQMTP3bQfG7j
ZjQRi4wtzWcJw0Hlbh+Z3xlfrnhRBJDdgbKV1PU2riEvci3kzMrpcpSav2+JfbjxD+CnVpecFE48
HpOw98b8Bat9QMGmrR7+jSqmCa6GXrpHHm1SkuaIm9M9UBtFL6eSkbG2aDrKsiFTpRaw9xV2cUfG
PRr5pbPMA+J/4HhrbITv+EzItjUS4zQqDdcxBkhlUdHjeUrrZ+XHka/bUjBoEzX1RoGjiWD9Kcr/
ykkEleUr5icKEp48xtwjxna8H4wfrfY0t/EQixiK0knPWSOSbTG/UMugRbpHnwRcmfWwW8WyqkuV
8yblmbnBdzEI4xmTNRAiNVn+K0tcgKPwX6eAvPxkhPgV38Wep1fN9EPHuDgOar7ofrpDNXCVM0Em
RtTw/dPdVL1osOjPyxlAMR/XwReWc4uqEqrunUrEUDOnJ7BMhZsBIOEpQBE/6pi9/lV1wMUQE24v
UpKDSQxuPEqW93szwsvSpc7Uh8lWqMxqCiIjGHcklW3/sI1qIq034oLUNDMhVrOBi7ZVJ3F/u9dt
d34oYaVPYmMlJdiGPSJkmxXFrcB+ee9R2BM19LGUoKPqQ2tGr/TVYkfJDJ1uRXTpeRhykiXG/1cg
0/nkMhKAQGuvuidMqbrkKd/BrBOdhkH4q5RNZR618jtmS3/TX8/dscE9sY5Z9FTX+XlupGuNsPIA
rK/i8I88ivoQRZKMYeQRVCO0xT3fNr6iH0a3v0L6FxFjDL9pMfBF/pvbokDjsMe89Cu3SFmH72Kq
Aw+kpCz4/BnXq1uZHqsVJDB7g3shlLjyh2HxnoC6774uEb85mEepnoGytLsP7zme+gQ/guH/4FtH
Cx35Iq9KzucgFrLmQ9VfiyZBOLc35UMIVvDlH8tR9MNzrqPlH7KbCPDAg5Hz8pV7dZeUroDIMeKL
Pf0LEpgKiyM3+nyvDjx85hWIU63EL/9bD1tpfQR0Xw1rhVkfoOSkPUAdwJZEoAh74qlRqaD1Vos7
wMG6x9rqM2zBDD1Mnl6UXGTMolPaURUH4nv5WW+Uy25t9jVyM4Dvesg6Lj9SZYuxzYk7tk9YC2bC
3rCTFGd1DwdwLcFhu1XFYVe5gc7ECpTkXoperyjYNNV21ZsADwzOBOlkpgfqgI7bgOWYgUJ/IiWB
5pmzByR5pKC8SMr0t6Vmhk/G29112+q6iKS5J0+REgXsUYc5qZg43TE6y+09uukdGO23XpLXlOaC
Tqd8krhoBBDy/PlkU9PURf8CSLAXfKUj8e8y7ySmgbFUbLCOtYkoiuUm8F+VG+kLEshgSpVxvPPx
juhaAiO/CJsQn2Xzw9JNOrBKZ5dAEtQVCo9uxdss3YWLRcAWgLKSd8NEn61h9vAPpREJIoA58zDt
3/jeImJHbTrlEQD0nzqWfcbys8lb0N4NnP40GIxiKi3L++eOR3jQwRaWgf8xHCuKK8TxoXl+GYpW
Tx29jkTPjBdSOAujJjaJqyPV5A58+JKTkKc5RVdIMz6UMrxkiTYMskOXVmRDnX5g0Xv0snBWTrzs
gVdvdDUiTPCZEmF25QtFUtW7qDOUQu86o7zX67cl0tteVLxbiqiCHIgg4iZbnqvkfmQdXn7EfATl
xzyI4woNwDOjAjVKhFU/P4z6grl6mzjgEQD+wRrHy8F5br8qfDyzb2M2WsP4o9jPxXNXxTir/RQ9
vU1cGuTIDwTMduLha/0g/Z7Y6YKOlNrVAvYp4hqG297WXjcyGwKUORr7FvTTwl8jHXKIlzmI1y6U
zTh4KLyci+hydwaxLwhKclbc5eFDtg00Upx4fvvXmSioov+lZ1OskaOomY7vb6I27efuTFowH5o+
/W0zT2u63M86vO5PzjJpTCuHzpkBcTTqEPpmPe18Joc9SEANE5efWPbgD2pcJS2Q/YZwwZBL2L6Q
OX1NbD8FxiLQ32fy5j47PRfDeQksAfRBtrxgXpP4yXUPaPBFeqV/q0bvWExwZ95F0D37ydPsaliq
su+PU3jl2ufK+aT0TTTicNZTdEs0CLZdWOiA2VqYc+mBuwnvGi6OGeTWJiCVb13ANzH9HOP3h9Vf
31ms5/9yDJm8Kli29WhbPhttWCaSgEquoXyLphZ3/U7k9QFbwvlxXl2vVHKyqJdNisLh1urrHzPu
2yez95oba3Ehm8VGSBUMerdRKROr4A124Ol39lyVrhCtdvQMyj1H0/XS4JeBDrYMqZ2qtNglmDva
/FbbRdCxUe/VNg6PjGa626e0JRWMZoNlTe52G4FX1svK3T4AzN6dXNv5R2gs8YdZcvI5DYIsC6n8
wchj2WtNhnXk3vG8ELR1rYbudQWV5Qrzno5a1xjWpIUDnn+tOAYq+ORJ3fE/PDFMinU+gYWpZP30
HEGi+RpvVml1Z6Ex11lGddb/dfwEreXkrp6pG8qNIQJNwR8vnZFSviCLKOlOimSfWp0DcvzLG6we
1hCGR7HlC4wsnBbG36p8iHUlTt/XnHyBt9wtBeY/uGcj5gRWUcfaKfrOmaYrCGci6P3c5Ya5gMVI
TYOp47rtkb2LSrRQX/SEX8PJT3b5TaYfDE7DAnYqXoeXZasLTCaxUC9bzIaJ3g9IaDywUyx0EPJa
XyylqBxBroSh1a6PQaOGefw/BHB+bIzBxe1XfKOribaLUTUqdFDHrR5iXXwAIcYuInUyty8Jud8y
SRSiALrXeQZEmi4QOBWvVnxvOGLBOvl9JVM3aSdMBNg+SLW1K9top2FvcGDe3194Dz08XMPU6Cww
VFdZ8Ved882wTj+KFVtBrcf2JdXacg0SvIttEsJGIxCl6a8TKTEjIX1EqQfJVSMcy4iXY9MPmWIf
wd8+vFUZ5txeaQhn4DAN00NaPAtqkBoNrGKLq4j1Ic2f7DT5MlS7yBhSPn6l3e01wmOUZURMp0fZ
Z/Rntuejb+QnVRh03pUM2lTOuddDk7i98Imyg8q371YdluNj6MwwbzyHaKGMGYbcLwlY39Vsj08u
zleCv0PgbjNENxHOUz0uyHfy9uBDProuKzGzmzyiTuwRA6f4Fllp39/DpbAhSC+GSaETZCZQpIa7
4CLfzXA/mrAxJAz9wNR8VC+EyTvAI5yKC64eNYiA6cQA0Cx+AnkyQAov6O42kYosBjLMPhiGc47h
HpyXUbuQwNSOXPJXVlloPMtAJ/1jewaExOPaildgQ1w2HlrVjArpZCRZeIkaA4A5RyH8WrHlkYi5
Ycq0I6OYreeWC957rLGkG0D3Wx2IhWz739HNEVls8kZGCTlk4esnvEFmAIgWMKBffyvkKP8hlcFt
QUsofYwLBjZrefiCflYiyqZ4pWRLCkkqLznQPC3inkEaxg+Ium5FbraY6evIwxFCLWob1hO0tRlV
+/5jEQdkPjmEJz6n9ZWeyhO6mmFTU6F+/5MmWdnQyClenT1haI4pQA0SgVKUSFPDN8P1ZaVFbzZN
1q///hGm+RTAXxp2idCTgSPBT6b2rK3RZpO1gjB3icitSp4yghrr8rxcJfgkQ13xvMiziqKML6f7
TulTo0PiFpgqt4bjJBEWYEj7wjUJkHsYMpASumk4GggnUHO5WBz79PFM52hhy4WQVkHlszS4lIkb
D9gEqVy2eDMgIM92mp0UpxHGdi3k3ThS5OXsoIdvJr6U3khIWb7J1GYXhtnis1IuDx6kBsllUG0t
SmQq2SsyXj8v2zymeKZAZaHAVgc8ZJXG0lqGcKf9jTAxkhW15VkbSQWWN+3pnMsPBt2gHYS4Ktk4
Yb+JiYw4u5PHvuOZ0gEpoRWMUSMgpYT+bDzWMWh9u4iGhsLg+1fdy9g639owcz6T3z6l4teyE73v
WYVzY4PF+SSyn/XGOvcXkcLzNBJEGGjQHU3zk0w0j3SIRRWurDSypiGDedg2u7NrFQO10mcXtWI2
HCFX3igOHC/xv+y1jUJ45dZC5dzQVltlH26EaaV87V3o0bn562vUD9rt5p0tTReujtaf5lqY2d2O
62TTjw/h6h8VwnZYmu+0OF1e7/fcRKz+VPr87TWHCk7k5OIbIuvCn/2llOCU1Oz9YF1svdJOlE6R
MFpXNkfIkdtXQyNTZ1nmF+zR37xyE2lpRG3BbhkxTnWkITnkp7LoS2S6kiqeV0b6z2wTQQeQSwgq
osYCicLzo0F4btCbP9ZQpQ9ZrRvE4tzD9W05Zchx9NpTxzxy1q5PUV3OyDWFOyclPzRbbygQhC7t
L3eOoOzympzuJqhDuKwh0rB2Q5mqISG2LyNS59pbZHgxgsJd+QoU3Pcdwtrzo3rQYBWXK7hwE7zl
qqfxZsvBLoSZK2JpZWzD6to73xwmVKzzXIWUYJtPAmNw4946cXq90iglrd6OWZfobwwxM8J5uzMY
oEUtJjOtHcUdoY0q66gUdM0NTRLtuxVf/r2fl1dedvl4WaFlqavrxaHc7l6UtVULNlkhIQAAIU8h
wXlXK5oGNC1dvi4BE8y7tD2ODQfbEK9vnfQdOUtn7Bf4tXZi57S9eGt8bO80N9tpI1MzRUSz8S9r
F4wU6p0J8seaARNESLLkGXHUtiE/vlfXehaJsiXWjUyoHwO2zw5PC8ircrX+IlNGtTKfxtJoxV9s
SgieD0Hfm0DppienTwILVPsUENay/WLT5APneLdANbGNdTXm5jqa8a9UHxwQ/9D5bKPXf8ZQF5ad
bLe8K7GzXxmX39GDAKi5G8u4ZSIVuVTonVNwudq2FL12qvlorMTXjMFZKc5niyk+1kIBfN6siJNl
AKxlM2cmIxfTKnTzwYZUchcTszLcYVa3ydbmipA4AA69IdIIzsxyKl7gUNNl8miKWrWfjKQGn3kq
1ziz7dGPWrot8n1ccrEM5HQ4PBLc8kPRYOVc8qC5pvw1gvlAaxkvNqWF3icT4gapwrq2x9Q3os8G
+sRrmCxlTaNiZWfzDUYMp5k6Zy6TBEayglFEhyIDBTzM/XA5X9l+WcNlcTqqz8+wj+LCuC4pjsZG
mkJ//+IYLDOFEeRyuvNORKPs+WM9PhkktPogKau4KXqfT5+Z+NCTooRQEi9pOTesmySQGQH0Wpsr
o5ibhPxpd0pU8kQC/XjJkLTHW+oZ7wBe26ECanMQCxqqRnqomZQ2dD4fc9K2fkYm8BCUnHUjr+qj
JnY0Q8ttWLyw6DbuENuVFb8DDKjSWoQNEqkYtwMl9WTJp5XhzYTPI7rEvDQQok0xz6X00XvMvnX7
jGr1TWp2BSZgRFP7VPE48z8fxJ8a8mhli4oHx38fQoNxQqsU4BYohQk4yF+TWNuW4nEvj4Jj6Am1
iJ/Qv05Z3TXFcO+IkeKeOXWrXKFlJv7+SpNo6K2Mx2+qzz5lFHczsB3sfXPdcbp6tYo7SEn3CBWN
rWFkPsbv1fo2SBn4IGoaF8y+OyRz2KEznLxYxiXb94ClFZ0DkPULXNZjccb5CqLy0H9lpxYdjBbV
uF13cttpKHWEeO213o9JMnPUeOj4IPpALGzhcnIcypuFta9ds+7d6EkEGvlHSFaQ1LKOJfumufwo
0gFqAjyRumq8Rjz9WEwrghfzAOtG+SomQ5WT9iFQoVxf8d629hwomxML+1OmRj5B2sHflxIVrsps
5UQkzpr/kVRrCJVKJG579WMmVASMzG+RMKeRpEJBk1ekgbVXqRdoqlNjajYxWimlOpybWHLatKwG
qTC/Pc7xwvAppY6ogDlw63zKp1qmAJYvE8SzpOHTFBYYmi2IaiWN2uYZ2VXTij8XZUIkfsRC6JWL
dZxjTf6+htTFt2AgCTFqZDZDaALAoihmizior+vqs2ge3V/alyFCQo3ZhH2uWP+yxevcVO6tRE4k
GGYWytQBfQcC6tEiw+eEZEPxWjxnU6BhS69GJsQ18e/VzI4mn3rfA6jc1Pfh1SrElfL6FsKcksmb
oxZXna7ylN9JlhxWVxmeIw9PDMBk1b4iIzWQ+Qe/vk9c7zOi8PkTEuj6V3ObziCw1bbH95eRGM18
AHu2lGUokzfSI5JAEykIqZkLzVLfcylLNnx6kW1RnZXV+KzcsmfKHsVHAReVX3MxmYmTLcWi8uoR
ElX7VGwpv0h/kLO9K3q2GcqT5X2croOJFn72XMmlvnWkXKhfJ2u1n93PGTfDaYWsiNaQ3vkqmerU
lXYShMT3GxmDv/FCSEb0F+tRWi2jQvpKUEVMX0fnXCSPYaiGMCZ73fKw3fu+vsqM+V8xeVuJR4Lr
MjyUptkUC4xCqoxSitEANWIqX6V8A8Eg8vxS7Y99sJDiyFxL6z+FcMKK5a3vWXxANIsH788ywuob
zpp2cbf49XTnyhILTa9Sbz6jjl7JfJ4+UCUh+qLJGVxAJMDvTWiGYwVx99Nyw9wf0XA6NiPsUkly
4PTGVRmP4EAyActZ7XlsfTUxHUBZtU7YBS7FcIJz3r4tOpX0vh7a8uhQzyfGXcRy7bE1F8ci5olC
gsbnxjrxf7nHf2x3fUB9H75vrWnpB58DB+EQHI2Voz9ufKPRgFJTpjREghztsGy/KkFIqY04PVWv
k6Ujv8SdTZt9rgwLc9XjfvET7r4MbH0B1b2AzAGLTAaYI/AhHq95gAbAqpPZ3qEs4Yb4MgNJ0jC+
EHQOUbmrLbCl/ewQaqRsv/9sQigqrZC49/rOpzkUWZBPqy8CA5QCWtNp1xhSprnFp5g/l4xHiUEu
QBrX0T+OUEfjao+mZSsBAYRp+yHV823+aFCoJCR0cjmQtqc+2N5fCJi6uMhVj65wy7peHsej0vMr
s5gniTozexFG6Cbu3VoJlr+rRTlCHN5NfZL2cwD1kzeUVI8A+y6v914FYfRPse+cDeodNT+76byT
AmAfP7gCYoAPCkyTU1rkZQLv0QBuclBOCrDp+uDou9U/Ap/XwZ17Ia30bRHdAH7mL6IVRyRNngjJ
ErH/71hSZ/f02HJXWjVjfrMZ5KF9W2eHgZ47GFfeRuT6Ey94KgFQS7PLFd0iGsAR2bgSTvFAVCU7
6fhjV6aGHKts9RPXerEUk37VIgq7g2uUCYsVYV3tNaWz2pcBwCJOMw1qqQpUf4Yf/Fzc3CSQZbJP
StcgvOw9ZG3hfJ5PXugSRakQgsIEOq8dQGpEu4Mxj4E3HeHyLGCEh6oYjiR/LxA+ZoKAUfp4w6Dj
BVu17KoeLs6iIJUDYqEw5pBgbDePwlLAR5cSm2hbSioPuYE7AbK8YAA++0TJaJUGP9Jauri5qf09
cdYxjTVTQhD3PI20zeRbWBG6yFnIAb7cgXDnEG4UYnDmohgs6ffnSYyCy5yhCay+kS/eREmDNapX
+zxLplauwhtO9AIw+7s/v3vYsHovhhvwBBVR0AuzShDBUm5v/Ugb0YCHG40tsghymqS0Jr8PIi+y
M9wWxyzZX2Hwp0gDvfz1+jtWNAIOOjXAy+9/EsJQ7oYWtbGwRamqH+rgnsiIlrZN2/JbavT+inYq
UOo6fi8uCNiD6yOZcbQba2L2K29cmwtVr8yFcvobZRjL30O9w+IS3KJ0cQU9zx3tMuL/4fzdoPDD
lJxQRaxFtXeK/890EfkblbGYkrUnRDzB9arhUvUZs6GGs4i8UCdBayv9zbxMTndtpratrcmzB23O
e2ixybRRd8kk+2+arUTdAvlhwotIvKoPL1mL2MCGWZ5dfjt6HAgcYSFuNMjjD1u4q0F5yEwFFE8B
RlMH3o2B4Q5NoBI5WMAVqx7VTVLueF+V4D71ivamFHdPTccU03reWtlAV0O9iqS/KAWyWLbohUJr
N/+EeEGZ57fdG4uNjCTFd53+rUodOo34NWvh6Vb851LNo6ZYrNwK7MPgjoeMZyGvTeFivnBKHMGi
r4q6mbfoY0ssT0AiR9M8umnUYxhYSNkoWoXf1EY/qnjgJJoHrFIV9Ej3H2XiPRz0BlWYHwiq8AEN
P8hPk95l3KbqONOSEwJ6opwxfq3ZnQoDa5NNhJuFlFYQrWGuYFUWGJNk+X3YamCDkLJ0JdR3GBoM
p3iMCXTmniRmAtr5nnVwkX8lP0E52xDrg01t0X749QPUeROxo3uvIaItr4XeZZ46YkSJXAYsY6E/
kT4CYjXyxx0X/C2eBrkMQyAuH8djMm9fJJ1IJPLUC4sCeEsPC/YImLns5N7AycRP0X8K7zArfYDw
Dw4FPbcgj0X3VAgGuknMEDWJiKGMSvBku0jxwPDsWIkX8EAwsXxt2AUr1omr9sdvxA/kRs62EOBm
zH6UVdeaFH8iYz3XdVk9FEICP18mC+EwNQUBeTnmVll9p4UXXgBDDp+ZgKEvo/H8V1J1qdvXktGm
Z/Ejs1v7HSLzxPv+rgQ6a4QdADiKjLKNdv7p6FaiTi3+7Lirbcq+U1/LjJSO7Jf1ob4f56I4YyWX
vj3grHwBHudd7ZA1JLjhM9hcN0OlCs7yMrSvul2s9RUBEOFYqSqtznwU3scx1HPbgCSFl6qtbCOS
3WlMl2/EpgRTMBTo0iCrH/92QMeJGBQTtXB/Dzh2rS4vlFBaNmuX/5p+FkRde205FFn1mzRRtk5f
UnTR9R6GTwITxahqK4b2zSR18NKSWs9YwtA4ZVZr6dVcl2vTWODtHc+9d0uRBcniDjOuNhSgixsr
VIj80BsiF+x3F4qzFXpHYs5Ni9tldrAySYhaQucHKTnp349mKV0qZUJ3ScN3BfuK/mvnMM+EKj2y
cK0SoYcme6otejMbisTXsjnV4G6MMI/RydiRz+s38KxkSBqoG58w8/zPN6pTRQv+VUcugzuTNVL/
YWNaHtpJx/m7UqFq19PXleObX7X8QSAm0qp1gtuChULVw0wwGmP5K/j8E2i6dOS0cjdf0adJqxY1
0/4r9bt+mXI38Rvz6rHtOcB5JhAL5d7cBW8TN5Eql75EMbiuYPTwYrcqBUr9M9eV58kb5bDaP1yr
L9Z6/oM7cfqsywqWoiOmPHZuutQlrYs+2l/Lfdlyaqg0TXvz7CgaJn/kRmiCTtDFAUatq9wiXu5D
/zCL7fmxhghNcNAmyzWnu1pDHDvCZYCdVRxa1DxoPvsZYNRtmGccNUXiOe9kPtKTD5Jv/+mmcFUx
eddWBivJteQg3Wnw2naUccAZgmFK1yB1dEeIcr1EqBbcZS+bXPMQXm4pB2YuW0T56BeTiNNayybU
Mg2qO4kz19ruz6CuK0wxGoJYNQojhMOqZKU0n3+nHGHi5hwRYZKg8ocZkMoDYBl8q0OveLVbRTfG
Q89oXC14kf+9clpxrKWEwxyGOyNzxZRuzpxT06Wfq/3Ik8r+fOZ0e/XLAj4BxzE/AWH7BnE6+Ai1
/2wP4Bz2z5iO9EH647h7F0D1DL8fJH+xKHpcUEmXxzvMkdffcye3w7Jq0QI/Sf/0mcPoIWfQc4Az
ahxjg12NzzDs5vB1LCoK6lF9GHRfC8PTDShg20sZxtc5pcIlnCwR1+iplHS1HLDSV0yPajqq6xg9
arZyMr7USx28JNjmFIhg3kxMZDsI6qH93WMk2fi7sbs1ge8aIXh9AHFC/dY8WYb8tGeehT3V7bZF
bwKH/6ecDQMykGCOy5ytbExeW/HYRnvZ30s5SPc68oHf0DnSc7yonGgBJrq3I+OBvjvB/PPEhe5K
E1qib1qZtD0PQdrNfpDZX/+7yWKw0clabfPK9p3VaTu3rdsjS+4cyUSuCN1zoO4jbGU2eTqCMkRs
3tGpNAID6O5McLa5G1BaziCMkin4QpsfOUSa92jiQMKcDRc3KqcHZvi5WcF030i0UDlbEzPrePai
mill4gcQ2QPs2ZZQHo5wAKD6/SK+KRTX2EsK2X4hahlqbHRI9pFkraa6V4j7QfgEIecL1M6yUax0
/QcUTA2jP24o8d1y0bd0eGRc96JyDYP3hpSmfZUOgnUrVfNq4J8yPV21omZEnj0t915UyY1IqKPo
BMp1mqpIb3ir8cIbztW1TndocIAl32vQlVihz/hUo11J2/FBVhTuggywkepBLqYkN/pPpjR3/xAt
c81kWfjNb2CAXJLILP62eInezjwI0siN39keugyRyDzbNVqbXNDQ3xmqEJIzZyxTlGfbKP62uJz2
kbRS77hnD+qDppobc9di7EAk7AIQNj8A7v4TIcTL0fOL6xxZ/+wwMon6jjB0BmvMegA6BkrHe+bV
pNWq7kdrqgH1q2GlQbdLmycmguWTNYFFhkmFY+PxXEDD8Ez4A9BhU++2miTE1mn/vdWwhsF6EdpL
XWTAB4A6eG/kNrsZkao0EQ4MqObv5YQnx7YlGmMlSM1ip/tRcwxm0w5I1gEjGYxHZ9o3oPQ4NMJh
piahiKEBpP5+hdWWmRRUDSQhBLb0pBh9zcNBZ/Tur/k4z4mvH5L7OXk1yPuhqvt3xYAHZ1vFeM81
5CH7FOa066R+nyTmpQlLDJ+4fVM0cwZVO7kSPGD28iVIuHl9UgebHstbmfOXUXk+YBHgfa4uJjNi
1FcUaUBgpzhz0fiM3qiUHK9Sffypy3/DUM7LT5w/3aOlfldkxlXSBTinYRREYIYxgk/HI8VDxLoK
qaRrJ/3qp5qDIM15dNup32ic7ythtuIiP2+E8vWms/W2DqQlIVQMWt3gnc+27ez66Yd2FYQDH4LZ
XRpDJYmMj7o01myh13TR3d8TGTRwSaSJ+iT3YDH90od18PExEUPY6dfAQoVLyGvq+fStgarmwuqM
+bU7jYOI5vzc55pRuOWbqHVgYypKQMmpsYnUPnsbTh8Yd4ODz2WAUtS0SbS3LiQpWwnZyXRHfRHN
y6AyGLzft6MCiBtVO+KipFy9ZnHCG2coG7rWJgpIx9llGO8G0qgdF9E0zEemU8vCByRm/RG4GW2H
uBha5rfI6lIMs0vvYdtYxYPLwXlbpumdNM4fULn8kNc0F7lERBmwe5QTlybSt6swfpFhUu4tZ7J2
mrECt2k7Xhs1Io35dfsbNJ3KUxCBMS9JMlGDrpKDyfPkqCI2XxITc4P+7cPg0B3VWF+YNMIAxLlx
4TmtmEFXi1eCR+LIOfrkY3w2nTgs8WuLKsojyc8eAIVfJncff1Gmd5gWKsDx6KMV2IMsy2VahJ8c
E2DVniClKd3FVh4Zy5trmnY40kNirZaF1XlZYOU43Rc/iqNJy678efYFAoK8js4BOsSGQE2UKwA6
8IgAlURdIL0m32o5UF4EAVdcS6g8CCWpueDQPme/po0PbFqH3uzSZdB9qrDyx5icXQe4FkUfHQnW
f9gPRzNsE1PI/7Ri1mfU9yrE+qSJYwWudq1X0HuVEejLw8OxrAzg+w+C0Vit3f2KyOD17ecqLcz4
o/tmUA6ujd2BomLrYF2p4UgSMqTUWnNDbS8wJAc+Xe61+j2y2uAy9ajB1v/dmiGv7Yj+xi8u2w5n
+nd+7yZii6DwsHLmBdA9BVVO9GwkXhucsLWqGyhYdkC6nKXmq11fChgfLusJaEbIYkB4WB2CYPtA
KEusN29eIhLzTqQlz57Rh5R5A2s5qdircR/Mguj7mTLWH9PRp8qgJLDCnVElu16MZg0ZPSJhWx8Z
KrYCy0NQtyK5K/mLMthT1OqhX76wb31hfMkixIGtL9P+sxXfBC0+CLhoXenUw/HYQTwrfrc6RBhM
nNK3xRCyT0T1TkBGtjFEiWybIFEaaXx4F9dVRdUg7MOaH0Yh+6NlfjR051krc57quDQcbeINhdF/
jleBhONSLg4jT2vK4gWiEsv2LKbSN02QidHtBLFKJRTnll2NZq8xv9Ugya/tyrPNjPPYBaTbwqLU
6PJIWt1F+SbPAtn6tNBK+iWqRQ1vKyqZYNyYMWL+eRjAgjr2f3y5AOZEGWRdiw4A9UvHn0FffjqJ
l/X79UoK5211fZlz1hJ5MAOrV5ft3M5OKfEJk5pFau6NvN6rEB4PJtGjlg2MhfAIewBGhIeVraYW
RHPuNLnLMcvTPVlin6dRk3ci3+RJyMKipOLaMyaG8AOY4UV6veh7ExhQIth6vdzGDavoIlIfIjMi
50Q0NLd1KV/5bDOcTbLe7PXEyDaIpvkR7F7zJParf2/3+H4qesKjDlFmxGcyk+7DLTcf1VN/alcZ
usw3IBv6hhf6fMF8iOjz423D0mwIKSxSZZcyjU76C/x0rt0crzmIkm14XKkcRqHT4ei9CJ6uj1vG
J7YGK5jqiLmvoHVh93AVTnzbJKkR7P+tFbcDri6lSh1CAq7yhotuQo7eHz+kIByJKHIcMBpV0PP4
S0SJYi5D0s26n4h630UtQrRafQYGcQ+hLJHENKpTMZ/K8B+AjVAEshCzjuyBeiomzTpku3tpDmcT
BfUISkKUrAC5/qbGJVRglzV3c6In2o5ji7rM2L7x1cLsm/w9ZoDolGgsCk900kVxyMcdiWnExktp
YLPukj2gUNlnROdwuywSQuXrUp2kGt8xuWq9q3+syuBnRsBEyZeEHMsU1Ilb2KBuTh0SnhdLnYA4
u46s0qvQ/zuguXXX3Dv/qD2ZrzpF8LClrAdijL8aY4kaF7zTlPvnKy3qwFaeK/fQZQksNkMHM8gZ
h7iPmBGKGav3bDXBnGi1Sugavd2tLxLwEEomJ8S7AzhTfsshAZ1OTSl68MfOqzlv8GKVJyTTeUKe
tQIlqE6a47buSb0NdFTZ3YEYB2/cGS1aN/WLmSFuVPXM+bEfZun+IoUQg9Wvh+XvgHQeOkJx/Nis
3604K9Rp99H2nbdGxQZq/H+B5+To1lsn67aR0gNviR8L7ZfEcWV+R15kVLWXcyCu1Jr4zJhmB1Jn
17m/WicFxyWlWo4ZzphHckIyJT/oeQctLRCOUFk/QbNVsfvwCOrmssXeGkdtFteF882+Ycc2FbSx
dc+NkhBYYA/n/+8pON27bnarswEIBi/sC+/I+hDKXwgAn/qPuA9G/EnXIerA3eUTrz/dD6+2AuYC
fsF26xDrqrvoCLHdueefyLYcYtUiGqAvej1Ja8i/xTJmrjqEdKejs2J+o/mYU4YXk0Yg3Uyy/CGw
fsDq89eup2zSyTTr/f0T6uPc+WfVQoN8U4XQ8cExIuzqwxjwFWQAcnld1qK3M4xNJhQ4UXxjT99C
05KJHpNAsYdQ6kP/hNDItv6psJbyOn/eMOy4B0vH9y3ZVmQdWrWOeXXm22uur9fiI2AlXnn7/SRu
c+WeMqZBQpiK+FUoIo8tVoI4znMwItiZVsciGqy/PI+RiDZ8DZdCvIS9dqKimg00XrmZ1XOzrw8m
ptRdP1mhx4JacAVXJJLAm4JhklnJe7w3zcLpEgcJqHo408T5jAm485QRJCIZiiRShd9ELGQoP26f
HXZPeqmyYl8b8oJ2/IMnsUqxVzUSEMX+C1urxH7njTXDaYG2Mk2w+xdYOnczD8tf3eL2UetZxySs
dfn9gKR3RVDqxcgb+BJ9qqIfeYK1GDmqiZ8Zkgi8Y0udxozgD7Uhm3BdWUvXMoG0x9DqySRwB1nK
ONAgNrI56AwC1kWkA64WAJ4rYJXGTUmh1VgiHPJTjZ2ByrhWzNX82hTiC6Kskr6DMXCJX5rkWt1Y
hSJwZkyqoRlGD7p+uQ1TBSEVp6X+DbkS/c/LoTSVCcFJszh8/rG+J8/fQWDmgGZdg6aF4w2FdFg5
weaogotogLeCjtvSMNHyZS9/uN4EqAlTEZ2GuhSivd6X9E4n/Vj4Gb2PfP8qAvctWlJ2af/LtWtH
GFckmXCtWwxCEk9L+fGDdiyoqKwfEYtNaFZy9QALlr6nFvUvkAy4sYdOzRM+p6+D2bzV8yTQBdFW
6LT6DXhe8fB8zK2z/nnajL7LD1xyMeNdSzfLHB3zgB7TN7izjsDu0blz+ED/S24GWCuLpvXQpkyc
L2kwW5TJs8AIv+l+dGUU9lavDG+GGISJGiZq145Q0lQfyRqacnR6DMNKU4COGKY6I2E6zrgngX2U
MX1KeF8AmZltxYxaLzDb0trXI5DeJurzzmyzO0MkN0ncaCK3aRVKtm6L5KbBY4cE+oEzNawOk2HA
bpvPJp++rbcQN/ukQG8O6XnOIkIca/qqydOV2Rh9gIbV7JCzpN+cdorrlF2qaVwg8zwhJGBqrSGh
ElhwOn8+lFsaKoiCWWYMREaHN8E0RKksHdqI3DjWCsxeCXkpAoq2IoAU0UhouqReJFf/keENlWLg
jelEr2foBxJCYhGzwqJe55INE1pw7qa1Sh3uNbUsN0rQxoyXsIKP+N/WjF/xF0uO6Nld5k9FWgX1
v+Jm7XUEuBEuIwVJMwNCORI6W4tZCfQz1OVivVWDjEr+W1r/wRMQFF/jg8u798ULAa/yjMVdtrTS
Pl6b8mzIe5oo8DDtogfuLruaxWC0M+kp1VflOrKO9mEQEO5UjcRXyAlFOzV3VsZ5PqqFU1MpjUVM
ydphQNCWFZWIsyZqIJgL79RlLGTgRBWWmprX8K890vLuNFHGLr+E/gfnV/QaU5DucPesMH4AMSEe
/UD0mrO0aLjqhuRtSPiL5FHz5QEMWZ82yrGKDfjZfOOFRaWmsDm/sLbm1JH0/nurHx1oUYJC/OtI
/FrtV/hGqDOv7+ocEa0/Znjyx6C3T/T6sIPthMlBBptVDkdSQpFQFK9xtkQyC1qJg9WoZqKlkzK/
nH48qG6tDWcInpFWbG9++INniaCUtM0M07C7u/+32qONlSGUZwgGgONHxz7XAEwB2ktuS61bZTI3
g7DxGVD1knOri5xn8inPA6687M9JwZSk5IERqF6R7Fr/CEe/p68Q0W5+oPnjEuS6kkL46Ummq/KQ
jI1f1+DpydeoPRPc0pju+RRMdt7ae5PKN1RfwMdMB/6N2Cv2H05Z+hydlC78GWZGMi8YKZJD7ihC
CyvYZJHHuYLY8dzKfoX+i49ZVhIqoSddrB1x62A1ROlUdtPa3L21TAIGJCMUjQaiC9ku2OqrhS08
agVG+/Jjsz1j1C6tkcVGB6FrS9DUIalBLRoGSDZpbpd+dm790/YejikSa8eAdMphqwCz3tOYQvn0
A9dkvzrQvTqleanWmP7xjmAbxcaUyasXo0eMyPqXMneOmzikYouooAnDzPaL1Bucv4umS8Ay2ZpW
fb9w4Xn+nJrWQTrvv2dTqNiP0xPL5h5LuoHjOTiZqFcTUOAiQDeWgAQEdCx1YpPNeZ60nQ6sqqTZ
5QnJdO1JSGtCzOG/zsuh7Yd3dWO6DKsR0u0MLA8C0SNhr4H4pPMYQkd5g2NikHuoqQ5R66Svnut2
EHjbk5kUUVG5xoN5W0xV66RxgiOdLes70HPyCBoyVXdWYZw6iQepNm6bukzjDuNWw1WAvxUX0ueW
0eeomoYiQEorc6YTtuoq3iad9SoRZ5DTLwkl/O3M8Un1fRHixZ+cI0IucVImyiCMpPNNxnCn4G4v
9aiSw6FTRecvqMF3m0SwZQLmxQ44bfD6R6sF05n8GJwlx7LoT9ha5FxYVhSpWkiN+caDg9wvvY5G
bKPx64/ljAhi3R5f65DmBUB85FnPtzX+iu7HQc0ciEt8EQ7/FlT0S90DfFjvoUQkckfNL1++UOhM
YdeqxvxWj2ZQ58F6Nz7ILP4MoN+rFZU8UoNS5Elf1riWyaZo+Zu/nu8OPpRDnrvZRVtBYGs3AXX3
yK45Rqh5hc0k5G589RvdRV0D4XXSaogAZp/PNWav8qYhZ8WRmXv8bHriv+Sq/l4xJYu2RTZr0Fvm
ce33cfEuma6auCImchDisrWsqUqhX+pc9OaoV12axAWqyaywCnOWZsLh5cjPTORoPl64wWkH+thb
iSIOUi1hkHAQ9zvVSSVQFPdRM2O0R29D8hz0JhHXZeqCIKA0pjAUR2b1An4O3jdE7PKBfZDRyfgH
VlaltF8qgHHqtSuQtwUqco3+OleVUZ9msSWf/NR/bQ478d4b3gKH8t2IPGGBY8RGb+FEf8G5kMaQ
cvld4G+BFpkVu4RfRdKzRGo2YVkls/FSUWpRGrjg6eYoxTT7YOcUEey8uqQlz6xTtmrxJ1wWE424
Qx4hgWZfeQmXg7JFQvQ99nusnkn63RR5BwPt+YM3mplG2hMKn2xmFXdsIatT99JRMOeVhrfqBJLD
Vb4p/hGVnfoPljA8TjzyucGdsaUDMrgPnMSdPWYcn/yl7rL07mnremVt9YdCzgECM4+DeoZVbxZ6
GVm7BnV36lxO6jfyVQxBAwTiVgDXV3RZ7KUKFvSo+4PD+IGhDYTtUzLymc0bM80easi6oT++0BBR
c6IBGQ2Hvwv/xFM3mS9VjFEGHuPtm/qal2fCjJBGqKyU3t/GPyOLkWDMBCWkeRfV6Z+2hdMfXhZn
2C79vQs6qHPHviSPkl8q6G7+o6cZjLca8In7zlBCOuK7VLAFEpN6w90w3Lp63XCkkzFwoZplFUKv
nnLdh6BQbpDr8iEQMKkIz/DfQY0UWKhcUCGCw7nSObO83aVRZWuCq3vdcGRT5uQcfuoDYg5hRYfF
t6qARV7QtxluTKk6zWFQ/BiHlobkem1TKKwCCfwaP2EiV7hmg74UgLRX5vkpoTXarxy7qkY0v3t+
2w71n/5ndK4skd7FmU+wSztp4g/kbK8lRZOqtJ1/nQn7MQ5W6Qy5lWkb2k3Vu2P4dbM6HOJNZD1s
y/tgff+SonIANx6v+vmkeYdqCVjnNGRHeo5hMnA/yhwajnBguOZf0Bp5zu0Bj6a0Ly/MckS6xnCx
1tkZHyOp5Xnr2Jy++Uw9yBIJvZBfSKwxhAAbBHjNb0TcVGj+X5+0NAsVdt+peuqf1YgB5rvaXQcM
difxMYylRDJlZ7r1+3Jv+Fgfh14HgYauU5Mju0Rul0uKVVs2AZ2fn2kE7uyvfOzzooHce9kJFC9s
RWDU/fM9is1Vg1pzFqjspStFHkOZe7720ccFCHoS+UdAYujkDnaDtn8/+N7h6x0Q9qWNzJKkUSGe
XEkWy2PO0Zn4S8ZZk6M15daMTw2KQUTbCd/Y4VxSEEKYdx4iscZ2TuC8vd2TdXHbWlTEiKFExIS/
cUBtp5Iu05L1MdI5eqbo3mm+Sc/QLiJsuxm5jALT9r2hOcwiGu3ehZgLwMOfwyIQSy95k/AApZz8
XSiODPKiZ5hgHb3uA8R8I7BohCsk56wPztQBsoO68h+iQGL3Wi/44BPUeF290Qf0uVAyEgRzgtuc
Ja4snMN9m4VLSJi2Yex+BfeHkadffJTx2SNDBTAtlY7rOIEWA40pu/whiEH2eAjLCyTyFvE5nUuR
CE+LROv8qM54UxddZDk7RJxungiKRj8MlZkKU2m78hbkdIWdknfZeuecV87mfQ1GTvOPTB7AOi/d
ome7ZqEfNXIPCmIOMHGLrEcUXdX1jEXed+tVJZBIqKvWWcsink0v6dQxb14GXUh0/goNkCfUm1wO
/dvlAPwy4Zo+Xa2uxOHDxfztPlBjCLcDPDxUXyN0EE+tbzy0LNRbLphTivfloKpC5rhodpBjas2g
LucBGyxbBuYqPhlRbC+a4KzDOZe60qsFq1vrKHN8lFL4sqz25hbf7FrH1rYLoFwkDqG2bMmghiZ+
N5Vo5Dl21SOY8z2Kh57XcBQtIv1LBFfjUAExHZht/wmy9rU7QQFx+R8Bagg6cv0Tz1ZiSvxnXHKs
+Z0OxTSc+qcdkgDxtDJBUHwhSydFV4GuCpxwpQEbm6OrWp0X4HUiBdTVi5XK6byfTBmpXzr480CY
ZeAt01guxh2/xHhGN4uZOvwern4E0KNsiZ0brAJS//doidTL+/KzCbiQ77dartDHQMlOlUfoPeno
GK/DQxSI6cxJ9iTwtlt5+1kaklF+Xj1lgcRM3c1TGk5l2E1xSMiTbAn+Bi9aSbNRkMySWbo5qJlJ
pBt3OGYtibR5HZWC2G/vssKhoVVHfAU0VbOxdRX1SyopAYW7StBxZfEuQJze8sVoyA1/9ipKZQfv
toDE/RRz2TFsxWcdDELr+Hkth/v/KjsmcHiUB92zi4e0Rbeuer3QFY8KenhWxvituH2pgi0DVCTv
TmIY5qNzrm7Xo1AWqhtVl+v9kPWbaTZ2m2jwxjcOZgNNcD0wmYQwG/I0oBmOr4SkPaN4B3XBqeoD
gKLDQhmdCkoKPH/ApEB/ALD6W/r3Syc+o6jwBdOTswGjQFd0tl7xpshnbXnHsAGK9hgToGKzfEk8
yE5YSu7sFLljQHmFBh9LUTtB4vh1zfcnXcYZGVz9CWiiW4Bb1sPXep5xcaGFlsYL0aCLv8PY+OCQ
bnez291JsVPouOb9+6wIkyQEmqvXRw3acJ/ew3H3/8tUlKweLexd3SR/nzvBx8HYb/PMEL7MvuM0
n0sV71xGMEZMfu/tysIGmqT1m6whHOOg/49kM63VqDx88iTV1rJHeGDhHOCkWxBhmYy4VdQWioBr
ujmAuM1yEmxOqb1MrLfLwkhTGchFM933VwaqbKavaSlPqfyLQ5aIFCJpK8a+v1gacOklJ6i0Ddve
pVvueRr+Vzlb+58kGtEcRQsysDRbT0gYeljgIZ52xozdojiRROb8YWgTTRwnyLwk58oNyDhai4wS
zUy8YPjLE4zvnAClVio5V18Af/TSbJUNkJYZzqUAVICOmc3QmLtD4URxZYNV52dvKv7gkF2QuYd5
l38j1Ng/tNR8kFRWpuLAKnWB+c/7OlW5cSSSf+kHMvI51jrmk01YXqBjQGMiB26RaM8niINXI+cz
PcdsafR/GjZTmmNanIVwSOhHvgHscsAuurxwMvO3ebVeB99JDZgfNgjf5H15OHv20zjFXhxTnlyK
wPaXYTfJ3fjoDNqiJECtRMGcsGQElIj9GeFGlWFXyO8d8TfzVV7VhMBcr/T3VAtGACZqTTFmPA8n
f2rs9RQbSS26enxcBW6LQoTZny/EBMPCbEHB6wfTPY99XSr/RjwgFIdEa9YHOk1Hf7Tjx9gYEU5K
0n6NZBqYxUq9NYOdzRUtMs6XCLF/l1X+VDrOBOW9+SA/ggriNrWJc0qGJSvoqF/A3rnYa5Jp15wZ
YWa7FcvgFxs5q1cz2SyrX128iOTEdkQUcgIK2/wqCGUcwVLzFFcpsRiyjbE6aM8jN4D4LcjkBml9
0wbll9sLiPCjWxi1KubOtVVcFJg+Dx+6bMAM9zBidvm3BvCkQ+ouS7DlERFcxxb1UwYFhdyB9ZbU
uKi7amzEACHH8yF9JNoF5Q055BjoEdynidZXpgDJfI/k0dYlbg7nhmB4qaL061SBgHikwmHCrKTt
lYeZPGOP1V1qKiKdYmK/l0Jk8JYWDA+EKWPmgVIJfCFiEjCYVy7o+NQeUH2Btl7AnuZ9Bmmt2+VQ
mZ5fIRvJ+DugfE3FlvATtgIR9ms5OXMHENNVIhT2tCQE8l5N5Q9OVaHcWN380+4+SfITGXD/37xg
fIAtTa3TR+qTjPcgaKL1K27SQuK/uasmTaMRMLQSO1PRnJyGAYpMsm2iAoH2P7eivnVuB4uZBVTx
lwu2l6T5brwKl0gnuONgjKZ6PCHLdo4NrtT6FCnhs9jSn6H1GJwQjenUGwwAiJtjlcXIsyJ9EZa/
KnKFi3qQYy7ZSW2BW5hNaWQ6q9xePE0XKOaf/eqiFfbMnLtioZB2QUlDUgCG+etTPpanc3xUlm4+
6kq+EhQGXSTvNFcGHom0EJtA2Ne/bJoF60RVZF3wSPBT72Bt0n/Q83mzgg77RjJKdmqbt6rOItBd
D4MhXTh6VuOqhhdrEVkucD/qrtJRvF9E9gAd+8fje9ARIsSEG4jIQVq5vWFlms3ijOwoOe3w65Cs
wiRTAmW9w9QPoy+rtfdFEWtJCa/Yko1qqZYVDO56enHspLKegSQJs3SfTdfW2aor/w4f/Cx+U99m
VuRu3+LxH+719wsqqSGRrQgR7hR3kLzDa0MM5biUlF22UThWXDNkVbrLz6/6bsQ0/V4ulY83c6Zd
fL1ilWJ8b+6z5+kSI6J3aKowIsUJsDAWc70gCVC4Q75sxCyJ3+wpxnCLB9/Jzia78efu2v5jPfRJ
VOl2fPs9ENpdXIKkFZgEnBf6+7mGlCwDzYZXte+JEs+10F4fcKuFeLlwTBqZ8klNqAKoer9muIR3
Pd0DOz9gYGoA42n59rXK6PT3c4qjYN3dqZwxa2WptvN6ZOUQX9OZxYpPVHqZ2brQn25I9800Yl9u
Lo/QvoRDbUmA6pqVO6bbMip9hoFKGzy/le1EoPSMru+IJI70/BkOzzAyPGsbgjL3qMgby5kLSUPv
QBxbX5e73etO30ZdVtmvDiuq/1vLWDN3p9z+lTTPnrlNMn4YvYItzXaHp2te/OrmuBBhPbH1SLKY
YR8c7jDcD5opqOuiMCkc467v24zkbgeLsxPMEgrnZklHpG+Jyzp2NEe2PVjIeghzhtfgS27v86zQ
AKzuG4mEJXt2ZpFC1PqzSOUbj/cqLPk1t4L90HuOkMtSq7cVvubw2qJudWQrb0xv56u0C7M0wVGq
9E713rkcbhFr5JwnS462IePz7bC2QEtp3OK39lWmV2g8XbR7smrZ1jnOSOrhEQ/wM9tkc81INZ//
b9N6jHXoAko/qhsYBqhawpVrZBW9zI0XlsgCSz+HuRptR90Emf//O8s9UoIBr5ehmr9OzZ878Kx8
XiNzCwNo+fx35BVk/FvyijYBIGsME57AXV33z1evVnK7QELzfODRvWNV7Qh1HIiMjYlBcPwLgRUL
MmnX368OyUAq6QpKMkIkFwfriGzEzjnhbbvTFS0+p4ukRbBtBhCXckKsg4LS4Z3txuRoywZBOUF8
sfsPe8Z+uRzgHaOP+A1+Lnb7GpofoWxg4dfgnU95yxp9yeCim8laTzZsOJcAXfC1XP6Xh+zwjVK1
tpmS9l5WQfkFaICJpDMKFeL2V4VUmImpY2dw+Z8HVJUz/3WLa+XHiYyqLVME8XgLpxqr9+uYr+Kn
zifSdc04gqfmSQGPwlMhEuad04sH/Zbz8c70zdMual09bweOQ3NnH3QkWGZzSEHZG5QoVlQGXxV8
g8lmWhklztY5yvJ/yg+y1pKwEJBmPvAZyJbPaIHOEyaJD4xExLKWjb60x/q3IvD1nv6e+Cp2djgW
r/qq347K8IZsOl+Ir9bdptSplVrfSYrup5WI7K9b6FVsWzfRLpwNfrS8ahSnPWik/uKnByh9qkP2
cRJhnFB9q5aNhgMgwv3+3UcAMg41Cze72n7QusYWcKZcBmZyTqUaX3xyKKIFhNgpivUgJsiCZEQZ
VSwjJX7NvLoI7aBh14sFnwBnwBFUYtW66BBulwRbHwz7m9RVp+/kmc1B8SQspBqCJ4PQm/Dtkpph
pdlS6rWMj6jVLSg/qx5tKdlq0x93+2ujOYUBprF7Ej0G9mN4+lQkd1rhhB/ydxxQVgXGdXYQhG03
fQ/dMjRM4djaYfS3jHhkEX0l/pWiPt2VXaROCJ+B1KXHURjLZVnzQMwSV3Q4MFjU7CdINmCfNcfT
izJ9MvVmuvLSf6qP1DFK/l+xhmH9XOAiS+jWDPNv1+KYkV+DgpCGVzJeW1/SOvkOLgf0HMJ7aSW0
hNo54eUdsQvkOV7I+7tDiQvWb3vZ/QwLGZkGDJ5em4SQfA/e7+gDVUhuj8RdG0xsVUab3y1TH3Wl
GpH5EdWhqtJRJcGYHJljTJsyPsvWsD2+fAelkkBWmrKPQ3pB+TuI2ggW6Gtpm9q7PVzrmqxUScLW
1j6xtsGQBwh0NUtlHU5sR8yAz9ET3JeOSreUK/FLBlccyCmCf2I3cLdbbrr0FL7u8m0yxwAKrMil
SqgiK0S3sVYp2ycpn+6dCPuP4ilbPyNJnLars0JVpM9dOxHQHNrwXZAo21+PWgd5qKPxQZ8bNf3Y
RuZ0LmBPpUQ+rLG39TtbA+6AwdeeMM008oc8l3bYFbD7LqGZZ/exJPgNAlaN6j9crq9b6m+8Aw4+
VbHRZpUEOPfeHFRFwO1eFj+qLWs9rfI9IjAR7M3gI3+NFyipjhuNcWFCuFeDsC8gUblRf3OtLeAL
dBGSvDugfHXCG7UD1EjPtn2jR09YStIkxwoGrHThVgNvxOlKuqmxvtU7aSm0HY73TwXfCUBEXf3G
QMRGBEDDZYUVamld9CYxsBcFoZX4MICvUt4+ClaoAhXJn5cy90SF9SCfP8pooqlOwydJGtINV0Zv
XBKgwZE1AKI/VHAXak882Wc77DI/fBtpTFeKgM8i83zOTylk2peOb/5xlh8nwnwchQZBCoVMpK6l
2kZkWJCKPQM37IRJtnTBj8Sty33CqmKQ2yafmTkLZNIXjIK0gTjreZ0jwpvvra3KJHeQDxNqIMCw
fQjXItopUf5o9yp1BAm2thiSrl8tVQYwuPhc/ksgmQK+wl+P8WEZkG7d8QwkLNTwObvEY5a2KTnz
F1qBfs5JO4Hy+3XLPPnEsbfrfon9TrIlPgbUxm2pVYGZgtvG5MKahMSKR4JmEVN/Qq+dgFtoroon
52Yp/6j3F35r2a5gKsXOSGuE/KUTdo4ImvbSiafUgSnpw7K5bwMaQSGLMXzxi36DRZYYQCZHqSuq
xhPD9pcpeNspIJ99vFBmiBHSKcv0nTut6MSaMgvN9Tvx0eheepT3BmWVGdVfVcRi7VeCQL4xHJIa
OazBq9M23tolVJRPm0hSDfWp+Lmq5AFc/tx23pQ6d+bfcBb0J7xjZSRg77JwwGcWp1ZDIct2kpdb
tUkIx5YxrTDC9mHDbyzK7tDWeiRYcID1b4Mxd6T3EqvnP+6Sq6qA69aw4QYkdB+wvTA=
`protect end_protected

